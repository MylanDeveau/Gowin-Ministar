--
--Written by GowinSynthesis
--Product Version "GowinSynthesis V1.9.8.05"
--Thu Jun 16 15:20:10 2022

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.8.05/IDE/ipcore/gowin_empu_gw1ns4/data/gowin_empu.v"
--file1 "\C:/Gowin/Gowin_V1.9.8.05/IDE/ipcore/gowin_empu_gw1ns4/data/gowin_empu_top.v"
`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
YJ5RXb5ESLoBVOFPUlewuNr9MgH+WQJfblrypkCBMyrpEP8km5PynWgnl4iG45gqUIjldOxD07sy
F5Li3LzuVYV+OKpZk7CZxtaJVhcYPHGD0CWT2QuqI+OYRwpYC2IxAhdNFO1o0/TOZSaYKDO0KTEe
W8KGgUW+RadsfvbTetN8BdOKlguqjuR3xNCJ5b92eUgqTUMeaeGD3jqVcgZQNPcbQ11P1G6Wd9yK
YvyCoekUa/ZxiUL5VPIzH6wu1z73fzbKefEUayYIX51Acd1ZQQ1Fe14/p87nb3TQRfo/T7ZRZ7hf
j/FlK31mwqUfnAGUA43va8XnVdt5ZASDJx3eCQ==

`protect encoding=(enctype="base64", line_length=76, bytes=84560)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
eMDMMdgUuupjiVRqNl019UkMB7eVAndA4S/oE81jdI077EhrWcJpYNoPR+PCayPoxGHxQgf297hy
UZvLz450ZSeigEAjeNPbvXFeJ+xK3B8p4gtcTJts8MiueX0LBcA2O3e7cnkUUrgSqUEsGHjIMVj3
RpCHMSo9zoyHrqRqunTtHv2YW9QQ0+jiMvwCVG/Oe2ofsdV7a9WHFlmwyFQ2RP0lMlz7GC8lUjd2
/pC5g/nixceyX/hLeTGhet7Xi2Ul+mD4EzE2eVQ9vWslaVe9VGYnfNVWlLVVSPJztjSucASUdS1p
xXevt5j2AB5g8DOPBEGCdtMZT5KaMUJVUGHFkyf67gfvLd6gqzMDObJcmoKytxiYc5OxBQ2/fHBh
ZIzvWcLmrgvTu9BO6qvKWQXSkhMVmVfvLDWiueeuXF9UTfjEixYi4t/2y/h2nwu9BqzzFHcbqnkp
Hsg1djUti1Gc4rpRAXBaduMEga0G1kxBcqxwa96l9FFDFOg7TyyTkAuhhgFpdrg797dLCrdIFz78
5lXRm9UeLcdU9UMXQvgvO4vWN7IyfsqhD77Qg84G6Itv0hhpwN6D88ZaRPg2+pZXvIhjzxKZkLpq
Uqtag1bDI33kr6+susUzxPj0KT2Avpr+4Zu2yCo/P92w/aWHyQ2YscLuc18obK4f4YxDaslPupEp
irEdrkejSgeIjL615rOS6GGRjtUUqXA/hCNk2cKMY+w8z9/309/YSK4LynfADuZKbLs7I5JzpE9s
g0vA4mrjrcrAq82KRpjQ6a2xqBfyjl77Ny84VUVws5AnxouaIyMMgx49IqhKQniNZLCSgNlenSrG
xREr9QAGsTC2/RURYEytd+++uqtMZvkCklXnSma/l/z1Vs+WYrkKbsVZwCIjhXc+aVVc3CLrwGKc
7HkaximCKmkHDFbtcxeW0VKwKU9Tcv4vdw63rQ/zq3ZJWmCz+MATnfiky7qky3fbtkOhiSDlQ6Dn
80wcfTCMAvNUfSvuB3qhIeHmVlQGoJ19Eh/XSgO3k/rqxXcEwCRFc1U/vJriQ/ZH59orsyH9xxrJ
ygtyZOGdMyzbr9s9nDrEyB93bfgHzi2UZbN6dNxobRXDoWhu0eZXWgGsGIoSTVvlEMDBMI1ANhUt
sE8JXm4E4E99evUpuS7Rr4+mIbFeUJhTm9X7sq6nV7cEKLpHggRTHH1/LTbmd1ZiGiKLSzOYIP8Z
OS01jp/e0Ccs9pFbn2FbXiIZLqXUniTtpS3lomfbAAzpyIk+1unsIL7/vGKc6G9Gv++3MQ3wqkyJ
xOk7axnrFzskO/On+xJqJVexfu2urUgPwuY8wIMxvw+8wvmfnHwWiCGyvsDkgj3xb0Blr8Hapb7O
McXTzS1QDPwdnhG/UBtIa/0GiQ8qovaveVmIzrFNkrnRqYNKnYsPjDy5hEsoPKxHiK5Hm06epXNh
zSDs7wdCvQVGgtXdqXZ0PAyP4fR2IdyU3I+/crxzTYJM6SbzaIAOQE9cOV34wAsMMjJu+va7oQVE
YbUi99ph5nyJCy5ZNsB6NjUO1y6X/S4dLDfq6kStJiXzRigH7S0PrHymuWx/xCz0m0gcebjcq/Xw
ljP5664gA+Nl3lGNT87wTkLrIKzfFKwLj9r4lkID5GhA7vx9oS1kgVrx8GFjq4rU1wZoObYDUALi
ZCq7iiVsWmZmh9wRJHvc3pIB5D7Fk/a4EbN6hU/fok0mwsnPrnoAZZ6/WMZmGl0JDJHPnJDJzOvM
ONM1ktpTVHYJ9gVdlpqJRVI1lWnTTcDtosmbP+95ciX/hKoS9jPJVLoT37i2BNDDoIIQFUbHwYPy
tZp2hpVwxvoD3y9Do5k6w2XvbwkDKns9sJjbGM8VH62aYUzF3dKdRNqsTck7XXeo7XjAunEKwOSm
MFmQ1oZZ5tYvbY7bhoVQAGYWywOfJ/hR4dhGZb4xuOjIUBWQ697HweXz5HayTevkfh1+MyS3SHYI
SeS6yosIimhJZjF250TCzhc7/wKlrNtLPb6nrjz0RgulxNFyvUiPDU2ZCw5CZxgHFWRP5Gg3vNVI
EMA/J7CA6Wmfoq2Dg+BcYApOvtRH2XU/L+SG//DKdkxGi6jRy7k3BvvJ30ul3USF7TYg48D7ovQ/
pFCvNtO4WcR4N0I/7EQPU/liWZ32Ki32iwwIatd9DxwTr3Gfee5vXDsAmxkYsZzl59x1CwZmjYKD
rgxkxtkm2eOoncG3+9VKfELz4/ePpdR5LAAQe0IOm4XNK0JheGJBXQbMRjXWrcXJhYdXJDX7REX6
kPU0U2JsPFJuYwDbBhwDN1icQYQC/GBDrH0m8WGk8+rDgEsvqXbeirVThUgIDk4+asSBfVLD2dO1
lr6ZrZ8FmqGME/UjarCMVmAO3KsajqHrd14z1l5BwhaB5SR0KIvvguXhTO3MpXg2nAVxKIlC7ius
NxdUxPOK9ij6HgLKRP7wYKXNiAoMjDNWrsxrvXFa9W32Gq3FddQqlDJWNxz4UwoNnYV1gD0GMmQ+
3MCtfAM4otvbfzuZC0FHHN1vt8huV8GOP3bKSFPp0MCDK/wilFB2xoB598kh8IgQmyaDgQbRxzxZ
UT2kbglvkyN/kSwwIZQLjUbqgPuRFBUNztfz5nGDQv0DzN1UBY8DP+CmoSps3yYSznVs1l+WNwzn
gnyydtR25iLW1kR5MPMcSZwewBVWkE7lnFK/g2HKSYVBAzrUlN3W9Z4JzfYo6vUkE6EmBWR9sTBq
paNIh1p9SbvXhutAihK88RHDLOtzfaGfVXtfCk2ivlP3MxhJewpXeGOcnWXVuXQB1mY52L9Fw88a
H74W4qlAhQjvwzigOOuEYSf7xzbtbooUEG4FFK/S3zyirBXmCuFHmkfaIAeLZx3IoRWMJE48qcDP
t3/+VBzIum/UeBj9FDOWJCpw6bfmLunShCsApRVcqFcnzASVEpuwH+n58FculAl2yHrUFCE7Ruov
OP5VqpYKOiF/RiOl7XdpeCC+5QhOPBee52Slm91kst2z2+UfqHYseQvC6xoOj7KLKKVRJBBrlwZK
BvFnkTrAPThpYbVVOSYEI9LQK9asqgtsz5wdhvE87ThyoH5mSxOJA730EuagXp5/H80wBvgBas34
n4YToKZ7vhvUD6HtE+X8mx5bSLnrl22sNASqgQkYRQqUzQ7AD/hdXHMDexRhjAx872WoKLc9IX1D
OdHUzmgwnBtcqCd1rOFEr3tPzKmqBFvNQvqkjoWrOWEcMEqIiaqZ+GiP7LvK3WmnQ6fUPQF8a+7k
dUBCIpyj0v5ywnABkUhGBjYMIGzjAnia5Q8iTSO/bNPiR8MuxQByT7TMZk/kT/QNjS4IcDkY5cyx
YSsXsBQNQyNHlka23OIh5zBTfdijpiIhkNJdV7ec2Rrt2zYfD8oqyFGcS3IB5am5KkoFk8p0DfEi
xjiAxrOPgCbUUQa+PYBdQkRyfKXHRVDFXW9yHMQLHBduNCFsWoL4xM2OHyQ5h66b47Yu0BPpj2Nl
LQlSoXYrdB3IHnkmMW4244ivZkKDS35UIkk54Nw5D73xFWQbXi+2/rnn3bkBbmmtQl/zL7rJtgbT
mMghHKjfi08AIxTo/C9lFG0h8RApjtdViL1heazrEQI5Dn8m4Q42F7WWX6R27UKDeNi3HitXzQeC
nznIFJt6BAujXRlELF0GKUT9c/JnH6eU7Ff78vorVF2vdaRgDnS2ySyZ0j1S+JglQgDGZRgJ/67g
2XZ9pIpv8s/0JkM0Fv4IbKexCF61FET480OqpOVotI6QHlMhIzeGpNm0a6XMwvzt3sYhRjaxN6fd
o05S6aN3ODrABqVqCusMsGC3GfI5FZwDB+WYTivxDUgVEkUKxDFWZWcVDWcRHUCt5IKlnacCSMM3
0GL7G5hisVYBV8Ut/zZk9zz6aqX+Zt3q14XL7AgfPYQR20L3nMa7/3hADscqJ2ieL0Toy/0xYxTq
Vfyin+Qu4Hp3Eak0FuBOU/+iAPRxHLGg1DWvFXDTQqvlW6V5DaiNk2omjTHoR+krnmqZ/+NBL0y3
Tq6C8uVJ4nY7muMbi7infmScA8ggV6n+IsUeIus9WepCxbI9KtuLVEBHJVA8tJLrlN+Oby7xY0Im
Dg2ujupIs5JUt36IuQX0EWcPnZb/SHMYq0Acpyld/0q4bbsmCv20xZUE3LyVWvuHRodwtWcXAoC6
Dsmqw/tfKGSzKs1zMQ88pxm+2PMUkxgmOrjpijz9sXvX54JiPG87oWSacNq9mERNGC/iyCV01WMz
cbofu4/HoILqD3XBgYKpt3/ToRygT9PsUT6ti1l83XgmmQLYvxdZ/PvD8vUXN7WrxcQUotrtRmUp
v5Az/CakejkzBqmfQfbMnt5Wv42n2F/SgzXmz+cknGH5KDXxyQPhGb+VS+clonYmY9uYT99EZfZ7
jA0vP7PeUjnn6+Vd0632f3nbaNchqdgY1GFxRQfFMAN/3Kh6gZco/znYw+co78j0RydLUUriIutT
+wSq1h6Rv6kwPUiwMInaas46x6r4ITH/x67bkveuPebA7ji1+dbXqls3sAlgSAtWHHSmmLbNcgjt
klz00gB2FdzwM7Z/q6JDSipNv+JOqlbXaS4unA/DcbxwbZ76VOB/sk6hsQeuwQ1vhdOTTfCGU6EU
8eeQhoNshelyUqxjqrc41iQqLwWECQhWtGj2XzXM4+X3Wv1rsWvFUXXfFyb+q/A125zVxYg+HpWN
xa0bwVHWtXZMTXylxLqNCeQ6AWYL8QffWPgHzOZu8CQx9ahwAu743FzvGplfslNB7YegSn1Mu4kO
V72ywbZP1gkyALHTEUXuwWy/0WqgBnOVUc32bWISWqAdidpdJXLAqiC/Z8WlTA6RsMXqrRQL2Jdg
S6WlHw+KcjOK18ZNtvOENlyW9fEqiWggj40zoZGmRY5JJ4D6Z8jtfMoGlv8L5+TEv8+R/hpNBk+y
oWQjA+asANFck4vCVF+fZ406NVQg0IrucGdgD8m7xAOooBA3NV6KMGzogB3/LYs9IZxyAwV0yz95
pnSmEF/UWVE4dALCs98EcUAKrNQm1rWMc12+Pmd6MSuFespQP4m5SIf15O95qL/muGa8wDnbHdfv
J1/OkMc0rLkbHcMzTHb93Cyzmq0poXEvnbmkD/HTiVXOAooBYPcggrQ1YmCelrje06LXIzRwJ+gK
Evu+uxkcFwYo/6BfMhikWQ0WQuVG6IP45seFuU3+OMnML0euQzVxcanPPG+As91dU3QAbp+tEk7r
EfOZXS6C6ec9j3ew7lLLG6+ES9a5aMXUVgiKDh0A0OVqrKNoJdnaYwfzAA1VszTmKac9Lw3Id2/U
EmDjwYHYWSaT+fgwciHGMtqPTqcV8qG0mf4ZwvtJY1O0yZoI3aIckfNxo4yN8WhSmntDFqCe5Fpm
NIFro3JQAQ9WAzLxqdbD0kJsPhuuerDJxj+kK3UomuBAt4EmLy83/ss7RLiDM25ZDLDDvv4nICda
PMKjeBsbVu/Xjy41RVtetKwEG+MZHjGHX63TVPIS3FhP0vo027OjRckRXcKRtvYv7IccJ1AJ6M7b
XPKbkVZ22JT9C8+lEIgeMM7k8LuyZrQAEqosClgpmvf5km4QktGlsmfENEd9Bn3Dz+GiL9hfMGsL
k5l+PSOapU6DWmtO8Fa7LFmvlzSl6cZ20VHTGoVkmZUrG7u7enwinAIuejjB1fWAj5wueWj/A4GH
iY4GyhQLXTipE/boLJddEXJoKiKiLwz1ZObE3PTqOMFZ6u6WOZRQJWbytOzzjTyHu82mXFn82X+0
3p8ROHMHaJ8ZYOxOUl3xgwtwsZdeWuxSlQMBYvO+MtVLRckbMsmkz+F8RGl5bCdBX7FKeCDGdb2k
X59EOj62pSVW7qbNZRh3kxMtdQEvezE5aIASSZ9GUsodGnKJIrQviQPoXgOuL6okdJlD8e1vU4Ou
DUiB5Fj6Jd8cHGifdvn1vtjNjNVu6YEEpa7aEMCN6agUZRVv5ffQpI7YsEuGD2uoxZb7dYZ0iL4d
1W5wv4luctDBRGC+WDE4EO7j1rDtdAbhUzmqfVIEpo1qpE/rXtpQfqFQfDN6VTAC6jJ6bHzgnTAD
cvyawTCw2hRh0QarIeakVT/f5r8c4B9GIn25H+s2Q23pVD0qGcSn9TCW1wHmDMd7uEPMz7HDVRVV
Y3cw33MM/bvUsTgzIAQzrg3zbNu7YzXdTIed2/HqXamyn6gZMHBayxbXApSTYZu+Kw5iQUUjYeH/
EuALsD9nUkh31h4SChTSB/K1211ZTdIc5mCTvPepXJ5qv5LMGt5zUOj/L2KTfT8AMKqs55hZEWPD
OdvCKnoZb0Ov1oAfBLxcAR3X8T7SO66+aV+Nj+UIo1w4mVeb7pkn5lCAtly3Q0s3wakBOjT/Fj8u
hxsLM6WVd0z3yGCCoLamvMR24MsdlrDpnH/UKib8POUEggft1fDYOQwbeI5wk6uGRX9zLIVZjZDG
SshQFEPb8q9BueUfrX3AO0BDccie47fsr6L3fs3Sj4bdn7u1NVvkvrfdX0NZV1GmbGTp3nJddSzK
iTlJWDRcoWavpmvVOuCo8jmNohHNz4fttImYOK04grK7hAucvS0fPAG7aXVf+z/x9EVGnqL01C0m
uEKA31Op3ipyJHmFxvDF5jbT84bxAgG0hHvMbwUpeIrnXVCfv4rYiWkSgcScsobOoab+/rT7CVDV
B/NuDiMdXzyBwjb3EGiblYlDhv+yXer6VtUJDdAQd+EJ67P7wXwEyASIrnnoGpGnNYEFnna+1hfK
LQX5fWt+gKkMZ8mMW15pHq/D1RQddnreGyQrHWsTeiHZQywDgdqXR3mzFcSlStTwvo9MVITTSVJU
oUL+ZtWcaJqsjqQQUKbGCKFVztjo69TEYdsukUjZE93vyjPvV+XqmpSqeffNAP/+EsQcXG7oOS2W
5DKCuOmoGexrKBbntd4IFkzlvC3ImG0v2bU8pDb4db9Oy4MUUMhVmuOAaMZVQ3bpcdGLjLYZTyJo
GRrjCNzcKObxo46IzCo0kcSZ/hyus7kZdK/0laEbBhumQvjJTRF8HDycNq5fyF+aOJkt1HQUCWzJ
/HcqGa7CFrKfWpA9I9g9sYnt6RtBS2CMHGBFiEm7997dMuzckHOFXnTjyzf6xbh9IwnJ/P7JSeeu
n7jUde+TKokDiXp1HTJ76C8Lb13yqI97zviFikRjTXVVx1EBbl+JwdVFQ9KAcOSpC3oM3XHo5L5Q
D9Af6i3aUVrSxwN1GCAgz9vvLTY93vo3zfeBEqCzVbG8gc8oLODmIsJiLDWWVNI/ZLUMe+z5RYoL
pYYckGEAzmb5igaKph1Z5eDnEfvoO74HxfEWjsM40lLC4xlOlW0GRD4Ad8yLmbnUbXkUS75mlEiz
1UcNOuzSTphH09UDO51AMDzCEWVMi4ddkUSlQG/aLY8+GbFkUCYZ2/yBKgo/jL7LSJvw1epU7XYy
zd1FTUsj6pGZp/w7YrAZdA0pRWdDiL9Pj669G5zvObvVW3SY7HuBaBkqTIb3z4hDRaO/BQ1E5dUF
hVFzTiE2Wy2TLQE3dU4hu/uLzeTxx+dyokKAvnDlg4eDIvXbAkqm/Qf0GDc5LxXgczBNyBtVNRzg
9pKcLcne3WW1yT+LUgnx5MNe7MGqSMt8ik7p5iHqjmt4yVk30SdVw6QAoWWf75IASnsdLFKQRWb0
RHJS9TXpFz45l8h3h2Buo8NTRa1C8zyMt+L89GJz0tFTVa5tbaz2jOutmAzLVFt3tNxGqlNHT2xx
jOcTWjbA8YFuX7FW7tmzNBM+eClR+qVLOYhbCderqb+MnlXxsuBwVJ6H9+yBFW625u4+FQumZnq3
hdSyBZYihfpesoFkUuwJ86C9ui8mdn46EAQ8UuEj9X/r/b+SjDulyHK0Ti9Bv1Umm9XaupJ6JlY3
yckMxUvKhzzuMZTfywbmpybv4+g6GKRUjLjgpdLre8pX7XI2xvpgUIBy+jVQ8F6dCFFuKVQ24ptY
YacKSiqgYxu6AmPAa9kJqxXT6Z/Z2iPEBdL23PQYOAG9cbWnEo++VF6POnRb67HRPcE5vXMEFwFY
Q4ZSEGt8qyFkzcaQez1L2/B3XVAm+PztSi21xRUnu+SrwkpvP0jIb2OhxTe2c7PuFwYHefYuy0dD
IzoLST9cjxvl+GBq1RKDld1SAnYJ7BJGGQcqVtIR1SI3bOdm6EICBda8dmwM06d3J8FRnni6Hx3o
Oqf2mIV4iAjNowUFu77uJ5cF0Z/Em6BFJi5ELNRt3v6nbRtQT0TfB2ITh1xo3mxjh1SDgb+Zlytj
2cOW5lg9/oLR3MzROdztXjuRuPbcaAgXe+DQSqpNXt5jRO1JKXbUf2uR4TAVmCf3Pr/H8+2F2LD5
prTQ0rfUMmbtigVMEG0yWGyz5Cp0btjLjRBAcNF5DuS/2viC1qC5XCDu2koyX/KszDPJcBvn+g7g
4Kyxin+sK9hg/43rbV6HjcbJkrSqs+EJGeajPxMO6xoPC2nEnWaE4U5POHZxpmODioETxwEETgXT
h69ymrslVWrXfZBqZVdfB1oIrPukRvCEY7lzIT8eJJ/ehAY0RF9ilfzY9eHeyt8+Jy3wIb4ISXa4
BkN87vmay5AE6PcaLE0U3RkeoDN7Ms57CH8zAbc6NQttgxOXQ1WZKHVlzR3plLrUEqERvn1a03Ka
Jk8R6BCijBClaCLOKvrnCvBz+yDXoB+zNUajxj+4pmZebqCe+QSPpzuVelfyZQN0hvuECUVRWgJE
VwVcDp9x7o0Wt5cRavPhoOb5gFHYp/kNapWUfNZqI+G9eyoPNdSozI2GPJGo4iE+azXKuunNfMFq
hBH3ftXcvFsQKZDCXN0KopLQ8WJjIilFK3753ScEf2pYjPDxWFdEIDA8VdGnqgDdn0sNnrLbEiUb
XPr+ONI57eoH1aEeblp+hGJ/RJ3jDs4fIlODrj0+jTU0bsPtXLWLtCH7X7KgKI4uiprB5zQXpwA7
MXw5jYsxns2J5ujVnnL7j/0pvoYRIAT52lSm9mjnU0Rzf3YjWig8Vr1OpIk2YriGZyBBuEYeOfC6
9J3l6ZPIuX5QZIXrtYtzyX4MLV2+23ZMyqYrichALZnn8UJMny+q+7IVzZdkrC9AlIUgoDmr1iP3
lDoGa9ZuwvhXdNKb7emQoS1jSwp5V0QT5VsSTEdmY9TX+KemCsak9Kmt5XI6Yyx38wcYNoN9OlTa
47LD28xwLgdi4Q3nlYv7wMpIQ1xugs0MyulVfjTQ0zBWq+OtmPGjSos9w98ZeSS7yec9vh7nuDMP
qxf0NREFBU8cuDPNvIM6hLm1tOinqDKoZEc9BZxYEN2RzJ1ojwi7YWM+nUMATnlZ+cX+kR2/bg+3
y/+mqu3iwng4Dzs3K5qAMViGvtmsyczWk659ILyevt98qLHUJYCXzJxOohX2GMh3ycgvIC/6NjO3
Pt37sN/V1Gp8E56pSniADiMcQrBo9stupwe+0D80uj7M901U4apna8fPpXMCnE4JkEplreCN3awW
IHHF6NGF7UUc/y/sJxr/RzTv/tzG8Rcwx5+OTgcFQsMi1sK5N1zWHuVq+0elhS3IPRJWvX6R4REp
rVUFlvhY9OxzqqQjA7m6Hmd7eWgZPDiUHcpI1VxOBe7d+6POv0rFiL2AiuKskpNySt5a1GlF+LFY
FWBRY1UIoxvwovneeRCj+hSH2YOx2F76UjlGjqk8aHW+tvNMudIs/5YL2wahUVm3hZdNUDowNW0c
HtLIIaenCIFWOs3hxO1srMA/EUyWDQ5ux0R4jci9/Yf00UhfCkQh2nDGhLiQ80w1936BKMgeSKOc
mqfMt+9sWdu2/nfsHsXUPQzeo3NTYcZ7GQQtnmIJoPkA+q8CgR2zt6nyU65u9kVQ+t+vPjNxNAeV
Ffz1i9+p9CpyZktiJzkzTczM2H59Oy5yy6M1dWTZqu6Qq7nkIkl4QBKJRWXEomTwaDwRNRX5eD51
kSjIRs6LoGaJpct5tmfcbhp2taudf8+GiqRUw8nDJBfdjVFsKF5slUNxRJMftzxFAh8w8TO6ya1f
w1hFwezwZJUpc7PblSg7ItHM6YQBzrJbbvmVCT+f+grGzrPdnXWUXz8EG59vO8bLxKrQb0aDS8ad
vM911KiyiN6fqzphijL6zifFsJ/fOYX7AonuP55j12slEbDVUve0sG7rdGOzuSUCPtAPPrnqpD4p
eC/LxeXbqkQDpgHIckbDFYr/rcrzHBVm/dWzCCDGVLF42+NMOmTTTIkz72WpSR+TEesQzWGT/bJM
/lJozVWUeAzqhZOzEvqx6iPiOuWsGNgoDTikVKukzpFOCK926BQecWVxyNnzl6JwDWZDsFMUnutQ
rMEbO1jIoizwRp97VxVyWYx+QWC2dOEbgnX883RE13aL0H4ENKun4FH6cSqAJ3KY/pDsKafzE+fG
Ksu/9lklyV5eYU8cEePitoToLXprbasphoWUHD50w2YeGF+643WhgV71Pc+R+zh9K5lRHkZ5UyZj
1dYyiUK7oiH376E31hsYJGauzPGZ9mdN25+/ObKfIGcpr9Rn+tQyCjz0LcQRjfPhlOD+PQukexQ1
NrTcORcPoAVROcR2fNpXOV3G3/UGBa4Tfk2ggYuowIbNy5gpCfn7/1SUz7xH92tQwSZnuqcjMe+8
AddaCpiwyGkN9GuKN9P7Aiu0ZQ1ujK1SDYGEidH6fBbVs5bKtIjqbHghvhDCKPXEONd9MIzv27fR
uOlRQyzmqvTz+XSLl62aroZq+6eN1GUqE4CmDk8M22CubmGTh42uDKEEvyTKgjhwvo15MkBmrnl9
htS/HZ9NoWt6PgpsphlDKzHm3Q+hwib7SOomBvOVcTtL+ddNYPY2vxNDpmiGye2W1zu0zR4hIKsh
t6jBZxg0oE85Wfp6f3i1Wf84eT4c/o0O0hMMcVkA1Vu400nr5pYF5wBkJqAtCDb/S7M0ulZy9q+j
NMQVIkCbFj+eZOYMJBavUySlEFZYEPqhR/YVf4aPiDTF1wvB1PG5RLoEv9vSL4M6UhC8x5OzE2PE
JVLV/ZnG58UU/Q1CP8VDa9QpD2nosQTsA9Tef89Dw5PX0cy6BBiu9RDDOszFSQRpTMnXPvwSW7ol
sQThZjT5cjz9PJeE7NzosKHtvYfKAgvxM5x0yzynEph9neQzNKe+k9+Z9rSo3xchK7wOs8VuQWMi
49ncJ16DfiFVFSlNcjLXlCXJepwcEcBuE5TdRxkph1bknVYKQEwdhratPS786184t9jWZCEWW1UZ
JvDSVvD1n4THToYU1myDpkcE7TlaGDfOh6UjL8O7gRpX9i3YCtcZCu7FA3QBKpt7S+c28vQmWdpn
KCZ8gAqrGjkuXMGu/ftQcX+Clo9pda2QT1Q41pLTmVvIqm0upefbT4Zw3XOZPHGqTJ/Ly8QMeyt1
vXn1gy3mFvo9Anx1P6VyZbuEddX5aC/mH7ZxSnKMI54Sd4sp1u31KmQqUB0nvHvfSuomzmm7zUdj
NgO7oidkRDgVKS4tR/c5Q4Xxlo3LCI2fy0EiWq/IGIMuX45PaoclYRJ5qCrYaZOXOt9jaKprslJU
WYfIh0HP6vDxlh/izwrUNh+7Tr7gNoaZx3m+pgEyqiY9QVvhDnoXycKMVr6X0pPMvhYrAfsqodOP
8BAsA53rAMtSTGUkPwGKVmwQWYcu4D2drtx8fJj6X3XVhtAiRpdYsSmZNyZu09784TNv4nVB30Rr
BPN68/SiROSH7RUa35DfPv1nzLgPfLlxjBVxQoZixWwjDno5r0ZUJ9vk4nBugjkHBwNoLk8Ldu+I
Mh1yVCrt/XVY8UDPjAi68oqQZsq2rcuWyPGuC8a+EAszldQYgyZuUysLjZidcNCMOEBkoibKzYx3
q8JkECeQuU5K1uIE67nuILOAykUzkYUh2le76LbTyOppfndBmldFi+u1m3QePJ9kMXPZsspCN5zg
VXuTIsBytXUoE6ZZDWWVgxF/F7qxrBapIQP18qHO+dF8fFycnsCmwss98ZRA5+in5e6Tb1On5DpK
wj8eg3R/PFxotaE+lauCnlGymLcjrHTWQCDJtdXRfoJK1E2jQJ0UIVvGxhyhKW1KueE5MD+Rx+Zn
fYGh17x+hFDO9YU/CMjIM8hK8//7QPVUhXsubuk+CdJMWfH41+rbwEHX983Jt9fYxcwckbYSOWjW
Rskf+Pv6gXbVv4gyx43yASwqSnx7spuYESKUH3BfWXCHlb9j7qxS9KyYmhbP9H8osLMdq7KvADmG
jSVG5RSob9s6Ymqh4PU9LIlZ6B4mHrKy5+SRBUj18io7znutaaa7qQBszZ3n+naQkp0Eac03cnax
rMEsxJCZIkuY7j/W76bX/XaNd8xKmRJ8QNhVF3BnryJuWLm8MlqThaw6JJMk47pHpRd/iOrn87+d
V9sxx4nGm0wvLTg3b3uaFkoeQZk7TAZqigwV4+TEjkftV1BYEqUla6P7pw9rxFKZHNNZUKH9yWk7
lenzguhYbqDTaWw50AUy2YjnKphDV/NDdAE5XYF+1z1kCFOV0mK9zIT/jThKvZxlY1xNDpXbJvUD
f2UlUVUiUug23QBkYjqQCOFKInNWnuEZKud7Q23kUw15MQxAUaHwZmNwn5odCoddvU0rK8mnbsSs
rYrBOL0X85/5zsxxjbaNBPTbalRKFKC7aRHTyPjVDlh7eu7tIlllLOl85MVpxequid2JsDlfFPcK
iwE/1jwQKcYlSGtNJcpTGp6axReTltdzP34ZGOkbISDcAC7bk1P9GqG3WXm9JkWhRs6rySolSOTD
LUNk9EL4qE7DUeSndae7pFeCZM5HoQOy0CUKWqpS0JFAXzHq61QfEpAOuCDVxU7jPDhHCffEIGZa
nth93Dmjm0bR7mZjAuF/IkrVuIEvhGjaoZH7VFnY8Thaj0sGUqeZ1rb84rVZZqIgx+3XJRqkUx6B
6P68mLyrvWIvP82StzxnmuA7Lt0HTW6PIqkuTr/oUConmpyGJ0KSVPOCjtpO5xPm9xQ8jn6kD89K
YtkVmsA8wGVfRgrCmTNORhzZd5e+0ehBHmDh41mk9/Tyq05BF6c9PLwbxoavR13qRQ1sYgGLf1wh
MXkOSLA7i9SbUG/Zu/+6owM2Ag6Zlv/Kxl/8+TN2J4HgTMZx96C96fUMTpjXppwWvKmn5qnsCG6+
z0An/ejespbZjz1Da6yZptBU4cL/NrjA219OT8ZSdWr/fV1MezBJ6cswCrtsCMe/zlIl/z2P3Bnl
IBTvq0TtVg8QQiHncHKM2hrTTo7JYZNl34y1dvBdCkyGRWcx0WeLblmWlk4sJpmMANqdNnfxj6VN
TUKP/DUcRBeSYCxnH1wEkO2N9S6tKD6s0VmXWfQ9+DbxjlMiV9lSjYCrXkFJCUK3L+cHTKYodfta
BZ09wpix58LSTMGhxKNMk6w7SVbCSbrZgCzrrKY9PIjpBgl07kAFiQlKW4KX/GLDA35i8j7Nhyox
7fbkCTa5tEGNp1H2k/pd0ZDvsUd7Hz+MSsShBUT+ax8xB0n1rdTp+M4EXcGBoVk7cQoyL8A/34Ry
6LfRoMtndVqoLcmgwrOiK4rrwNxYwzz0oK38IXkbBqELzluIXIAB031pr4j2RBQeDIc6mMt+Av2G
657e2uetkrCDy7iAI1R/NwZ/N0Z5IRsA7xDOvtKJRGzlxc9tEFnST+Ny1gSB2+/SjK2AbwABTyd3
6OxsfkOgjEs3X3AcdwTNr8JgsGyEcXQhijtBr1nlXpdzwA5JPOjHOTM4oJYPPzimXShWkpyVF12L
/6rW4eY+a0MD+2xVpch8E4gwLyybLmhx3KDO+fMnmPJ/7nsRZpd7ryJDkYuzIjEiHHQVdI5d3VcZ
o3G22kqUmY538AxZ0pfJuqRZX9M2+AELWKUM2He/jH7QN6QCtImC1HxS4ziSuyrl0VUszQ/rjVzq
l6F8rsWyw8vw7eWy88r8HXng6o82j8tRqVb8tf9FWo3JRYR0roc793L/eLmZW8E5lgmmHzRgG0fW
m0DrMQmvTQkbMDS4XI043OoR2Tv0DRt2NRZvKRvhx4Tb1lRhJNUkULxO0qXf3/JAhg6HH5ZxOqYo
ili44YmCckAqeovLqb4o0YVLBLlm3Kj7BpNh5J0wLx5knvQ9YfZpOsrOjSQBJokFqc+Cep2wZhHB
ZrGQPgS5GVrb+Adtiue4ycPnkMLrQmbX2vhQJ13Xq0sBzojlS5DoNpaS061zmh2P24FuUPRZlhQr
d+MLFd7FwqSyDi1sI5DazcMY2sjFd/fO/3DsX2iW4MIhic9Bj9U8rM2YfsQvK2gMoaiszFvipcY3
GbgG8b/6HCKaXQQCEfenllI5LWNy1kOJgyfLkTgsVCAA+Z1My3MeSnucMh1Sd0h0Aea/srMkbdNC
9Wco/SuCPx8pnbdV+gLeR6NNQfhu3h+miW32VZXyILK2/jIKfx9TfjyeCP9pk45g5kVu4ynKQ0gY
eT9Afink9SvlIgO5pZMnkRx5hVJ5UrUXruQ5bfG7yxJ+raguy0ASvjsOh1fvCh6ILjqPrMTNn+uU
xYm5ZkpGL0rZeaRKHbwJiDjYOPnJ5d1Jnmti7QmJrc6rWu36wiyULhjYVUm6LXGvNhjtH6bcSTu2
XJF2APqK1BqOGk0w7ZdkLwB1myq0zwWo7oafZD/fRDR7qp2/zwELeC5//tHeeTXJ7UXGfg09MQto
Mp+/db7UhPu+x6FZEbhUtp3BhOqM7MdaZ9k9HjekSRvELhLnFpb7rXJ6aXsRdzO3XiF8vVQIhAmR
7jNhkUC1dJxiUJj0buUts2uPZxL8A5mGHJV5QMaYEhSeKItCPFzgXxqGdSb8R40ye9wbZ0QGcxYT
vhtQKMGOS8kk6ERRqse9mrX1+Y1UyJuOlgdDtojUjXfnWxMQqdFMnVrc9BvrZvo6qvqvN7fshoWl
VCEIAmTvGkGSUyHOWnmLqLMrcRLOMX1u7t0N628aLv/UvoQ7sPWYw8h0OhCpgSb1BztWIP4p1VO7
lr44kEIlkQKFLvXLrCvLEzV7Ix+Ea2Jd7iMfDLrSAKQO0WJ4HGPALvEfhXv+sixarVo7zBN0vp3E
74fslWr7rdTKaouNkBsC4tSEPLILSVhoBaD5mxkybITfEbAxw4VdJHvsuR12pXfyFquZM0fYi8qb
XONoMbw+Toir68o/4QT34rP5SRC7UmS20J9Ls+vdx6X0xcLVUjUecjFJMrUwUC+XEL16ySS3Yg79
zYgXwMUfPtPcHV5ixBKl9s1cjUrmkeNglAaTehj4LCMk+wYS42bohD57TmCGTxyFZZpqRiY7rb4P
Ia4rG9R/zq5TSQ1lE04lHouWAbQfNPPDx1o9T7V1VlnUxyUzw1aI76w6WhOt/yhDfWGm+ooKszE4
jj2GRh3LlZru3YvXy5j1ABNIH8v9hy8eisPnHffJSbDhFs1pa/HeMCDLmSdvdQezhbj5eoDi72Q2
nDfX4ANRSTvIr1+pemSsYH862a4GG32X3z61rCrUpjys1Gebx2sVVIgoHah36Tf0vA2e0p7OQMgj
A4gpiI7wuaQ6PdYQ87qEcvOIW83wOmF+y3nwH75RNahUU+1+8gBnFlU2RFtfehQZtfAP0bpPHNPU
DPcI6H/AM9s41BUFloqkfZEWsnMrHlV6ZxJYiYNgzuBiiA3OEL6rxA5q0W1k5IcNHAJHZ7B/kxLK
RZb8oiKSh8lSW7pycppzAtDyYOLhy5EKKxmB3lI0eJqIsOqU0Ld0M9TTauHV8aLYtATmi5KOFcgD
VpQfHVHr3bQtuxLLTL4oqDMXRViljn7eTsKkfc2Z+fneCjunQZHEMCU0Dd7JnD90zXmudz9eDeL8
6s8YdkBoAxuOuka/1OeMvOoSObSh2xC8EAUmgRHIdkmTD61UkwieAUdciJTrQxm2wk/Um0wJySsu
+J3IYB7V8hTmMo/q0UoGjQypOkRX0aw+KpYxVy1KILuom1IkBBV7vlOvsePefCe5HWSXfnY2C1Y3
fSAmfKrJJ6oObQlo6Px/DzkgAT6JRY4cCXU4EIQVLpyulDxUs2ggWAAcmpEhc8cgfxzSIi3/cQTy
wr0x6CEFyQ6PBNbdhtzYr3hF03VbTNNsvzst0Up3leuvrlEhUh5WbO/5bIN4m6GHGmu+q7iPej9t
zr4i2M3tSqA6liAZM9BK1aA4j0Zi2hE7mbTSTdFnIRhxnzWZ6sD6oK3t7RZYHZdweu1ESQsaNewr
M9A1NW4phiA08JnwKxZ0IbcRnxHIp59jp480DAJPditO0cjQxe/I6dnBK6US4HnxJ8m0hy4KUpog
uZpf8XUZfYG59Dz88QRsh5tuzzKb7mUHX0Z+FwPvzJaUir1V+KD0Pg7QQtmronzf3wNxRo9oPoQF
nzyLfWM8ARChpaMbZuhtGE4RORuBTdARXg2g2glBhD5XBArIc0cYmp3R5sD5C3GHb/6o/oco2bgz
Cng5h6iC8kzh/tj435ia+jrihR/sB4/wNB7jeWETouP9D0DHTwR/i8pguqqz9u35wQpRpm9u9Eqp
jCYXWqhkfpMxMR3o5KuJPZblCuarQoGQxgh7HIo9gb3ox6bLHcYE71Acz837vAl3nmUIyf7yKCLT
u9Hnnsz9kdVHC4Kc+fddPHCTx2PJy90Nc4o3aYMKPkxSW3aVQyX44EZ35VFsV9payuNicPB6GFAq
q3nMHxuuxYWPSVSWQp6ij17Cfu7W3yUfonxEeqXmkwLKPQ2hQsYqmXy12tQr8CwOD8U/dGGjhw7o
SgEwEmfBFyBazaW8QnBO2g4TfX11znXuq2QgPBsVSvXmB6XLk+ErpphHqYmO8X58TqAN000M9ObX
zE6TZoE/9AzQB0MIiHsOiDGqEoqvPlny4cx9cAU7KRlM94eV9QLoJDz3pQV9USqhjKPd6tc/maYG
aCgZnnGAPCPYjXPZHhJwWJP8kLBqKLGDUocJl4yDc0rii03JHvNYt4fr+HX17wq1AgQmh6ws65h5
2XdgykP5sXSxj+3W9g393S1MaClohexTMzsIRS85rhEdhjLk0gxfiUO62mCrG25JOedFLNgtF6Oa
oWFQc6NS9fgEVfnJDL/Da4kkntSf1wuqSsjcKTDMqlWyve5GDr5gdmrieED12H8GEex37uS/HCq7
xYplu7QgQLGZkxrFp60DTsUZpt4s3SyhllU0zF26VJp0sZNPdCJ5vppDzqHJ3xc2BfbQT2lG1VJd
QhmtE+CH30ekzfQB7Sepzj1kdPgwaBOZGEPGyiD1wYhFcYhd5cS48kwaRbBiUnw3na5jq/EZOmT3
bkyHATJk6TS2uNWbXhvJvlIfk0NeL5uOI2JK5KDSo64RF5RvHD1ewMq1X0Na+pmXjLnqANixxSQv
jG8wChNRp5edtBnDWvMa0mP1zrNTCxXXaH4ouSWxVr5LaJQcW8mTuHcUHIFrDWFcEwFlDpQ72+n6
SHPKiGYs+8iFXjJFTmGU8PsqjRWSwiabzbzZ1vDVaEC7rrKMohYHBEm1oN05b0dV7SeumGLtN5GU
fyN81BqCE9qZsdkbsFHSfVohhJHuMKS+txuE30lhePYFsCfKrUwcdrN9aCRpcq5qiRnGwzwNjypD
UwjkFlD65u95no540k9vU3iZlmQOCLpuy/XMlBJk1rvJ1tS13iy4g72cK3+Bmt5vU3KYqigrEcZF
zrSqf+xWYpHT8Ucpt7pEAYvHrp0K5cyotht1a5o6HsnovJilLREjLoJp7IF0r7PJZasuIsCseJH8
OEuDgnAFD6smInEb2qL/a7S2lIRFXJshf5zlr2KfzxrJvzl38F0kErGA7zs5w0gPmOn3pLqRqdaS
4u4JzseK4U7OhesewpDV9au+1TwhAXqoC6U7FASftNkm3U8B9XOxEmt2aNhzxUqWmeMEC0QhO/LZ
HyVF7cVFs+63bQY40DJz1r3NzdElRw9sUWHVoQTHLSbSR2/ZEvZrjrK/fe7qPPfwO4JQTKWH2e8n
V6wirUAYDtGg5CsVevGPQonB3DYKQaRod/SYTSNcf3HjFn6UEg+KdHRMfvQM54r3USrTJhI2oGuj
7lmiSAIhGIYNqJ0FBBx08UaZKaW/xsDhsp5kJqpKss4I7RXDF+d3jGgIXO8Rbf7xQoY9YMacJzpd
X2cJZco0E2625CRaPkZs+ucd+jUp8bQkpjKan5SE0Xi5ZetvLMCabJJJd+bmHKC8JAXRI39Z2VDY
yvwFXXExBzKgYdAvyo+L3Bl+mEIuXGoJ0L0nWK5MBFUF5QT7yQr42wEBiekqhiAAOfc3+Bs6duTm
6RLPsNeuSnGpDIJuuQa6qg/SQ4pSzg26FwHfZYtXLFpylbWsbsU6FwMcCj0U6V4FOFLw4+IJyIur
nAOmi/R82waWyGIAL5r6JO+wC8O/9gfGjfH91MRzNbl910JjTU5XLK6ND74Vnb7vd92uvy10EsZm
Q4QC/DZzhMRe9d6tNXG+ITFr+oUYeqiHc24Xf6Mf9vOMAt1n9pn4s1fHtTj/fbl/ZkXjEVQFm58J
SRu16k3UDBU3T7I43RbtcKhv1K+yMlLatCrCdKVXyz2fJ7bYRZAC8FeYY6MTsQ9YkDOMgUhesyee
mnYHhQwHvdOHDp0TB67MB1pcuxffCYpWWaKA9j6IAMlLMf9742zY7jonJKfhvId+7TMKOs9ID00p
Bo8gzBxluGIprgi0gwykx0V3s9Bd0J4XB0mHOD6rON/bqw+VU0BUzWSKghZrCtMvbSaDvsZPzFrN
nv0nV8QV9mORKxNBxpwRNnFnzrIUZ0hy/u3UeIZ/AxaqxFPU7SxvxQRFyvMa3kUCYAcDhogzb1dY
aMHk9ddBvN2ODjUeY13gzXecjw7pYVVesishfQdc+6G4HllxboQprDS6KUNGmhIwUGbJKXR75aQV
tMvYe9+coIKxrfki0qcdnI3lW81H1l4ezd7a7gNQDcEGL6TaDeqgDJIEgigS+w2jOhRWDJPPS3e4
kcQo3RWU3cujRXew/D+YyMBEbii5zOvPzkBZAal8HryqenMRc8tN3MVA5J+jxgrSTufm3wr2zXmt
VU7FcVhqukYcw5O88/JomKZQmrwn6urh2rS8OC27f7nDvtpUZnyxvX++rTCu7KoOyCoCAK9Itu/m
bJf9HEYWg1DYl3WwnV2L/T/rTKgR7TSPc0xP24qKA3j1/J2uWLdilSi2UsLV8C+1m37SmZBhgg4W
GFTxSSn7JKtBdSzho8mxRARYWeZh+VDKb2460Y+UicgLdG77KcL0lt3ZVjvn4q1pe9rzCimrIfnR
lTqnTZfAJkxJBawzwr5bbXJ6jN3ozyMC3Hi3bl/DwQkC7CStb/y5LdCCaC0kel9uog9Tz5DQqT75
WVHawqZMiAF9VyIscN1ayIdKYNpnQLzxDji2vhxN/6uAapOvtIbh32Ay0tiDjOrhVh3dNoOD9Gob
k5MA31T/Cv42WP5paMLs5ZURhCJEniKTXv+qxBZsG7k/Fiy9jekLcqkBUgSY8APtdnY49amQ3xEj
pGosGK2KSWtH+Ua46y17XF4gbLCeH7KsuiDbPb7Oned9SpXKvbdjhsjT1PrBag81ONHcx22IKCJn
VLsJsnqiT8FfrW6n9eQgExnQ1b/olxhy6MKlLq5IliNuDHNRWjDL0JCk+Ne9V08r52SJSEJWCxwv
nx3YJnfKwFHtDb1hbTuHkjNr0/cemD35TqtoifT9O3Swi3G1vzYvAiD/6Ckbra8LI+AiDtHdadIj
qCDji633X6Su0Wvgf7w1ExcwJK+YJohlxdVrBMsn7jzQKibMvqy3In0dUvV3vDif0dsB6EXXY8I2
Nn3/pgxAwNaEZi556YQoSPQ3IOs/tNBehGIQJUUhosdzD8NKHFfJCuz82sAJQYui6TCtcfIUndU/
vu0cajKWvesshZpXhgvE1lOLkFyszWbVeXgGqWUO7l5GHKBS7M6T1Fy8Juk+D7OhDpG5apCpL9sg
S2SuX0J7kOFHc2hPoRu6g63otmMr6ybsBKeKtlN5pfPlloznkPlR+Gv71b414IBo3GJXIaH4ZkRz
qgf/U0sxa9yyY1p7GXf7l9erFr9DoGbZyc6ISmKUUVCdR22HC0o8RVN2GXhVsUngO6YMvExb/W28
4SnlJia6jUoU86d50o5CYjX0n2r3G2j28ftSWbxjj3xMV3vQC0FPOTrK7R84MW0KP2Vw7DHQHvzB
SMfCMqZKDoBQsG/fLu2hqfbDnrDwi+1Y+NrWfhnFUCoP1Z/aarD5c7XQdz7RU75qhRxjpJ1lpgd9
ephOA0uZQz91At0nUwhRoyqOSx1ir5uV9JrfRHsHGT8gu/7Vsv4WJ4WPDfIh+QoM8uWyZkUUohKM
fBGbpbEh1Q99Uc1TDLxWjQiiZnlUVt8ZtiRim7XEmomq4EqN7X6JKlagpm1F5Ds6R2qlukGXIDvL
MBOeR1aXwDIHCKpuTBkV88dthQ+F0604SeYHkHQwtk9QrujBnaNlNZq1VTUe5oui7gtPOEFiJ0tr
QSfNLvKgs/ULUityWzm2aa3m0xnJeZFnOPO5KGAGRD9T2oG0zsOtWYdtG8S+8CMZsxlt/9Ff0KpT
nuvptA2DiYJRbK7NkuNCXbuyP0kxc5G8/OeUikszs6btRIAeU/4p+PKHrvchPmUkhyr/B2THLbXf
XxLvq9j4Pl/2n+UaqjIY2O9zb8lGlGJx1NWXAr8J+JNSZvbvcVkz4QkSzesZFUjRdgwXoYWM5Oq9
TCvDGPUSwmcDGs1BPiNy28v2dBTfVZTRETyy6uPgkiTppP7xj+d/QNL2unbJrseQ8tg/8cAqf27z
LC/fXkneAd5UYk3Be7Ea9ftC/Ew3TvE7ih7Ar5XCjvLVzb+2uPddSoXVGH4f6HR47AEq9AjDOA+R
jq7t2FN69z7kTxJpB/1ddE2pETybd9l0wPV2yDs3b2YtIs0CiB6+lxLfyLTgBtjLHlC0hsJMYH+e
QiYgGrD86d7LHRa910J0ha/fu5AuEttHQZ31NMZ9sMREtlykIS6s4g7aCknxoJ3WBdCQ9nNNa0/B
oGOJ0Q9vRA2Ak0miN912qOz0QGE36xkD304xFV49XWgWZMirB01fm5n9TZK1n5Yux2OezwwkRoPE
YS8ATGMftj65gGbFHlVQXR5Hnl0119GexA+K4ZIhZg/ECPMSFSPl7Xj/eZ9ivIryIELvpMEP89Jr
g9DsdZaSc7p6X0XadRWnnAELgCSMfPhvyMYEmllQRA8/DSr6cL7SkqQOFReaTssE1C/z7vFZBq0t
nbHvDgitaVCYz4S4IJeek9GyADhO+UKdFlIWeRt8jetRS9uo5M84s6S5r8lmYXQ+ZY2dP7MSZALx
baH08C1iBfOT1MWLkisd1egYPqsKEk4PMvq/+RbvPdvtBNnn2WhfLtSop+I4RsILI8HrmL4y8XZo
zPrg1dohF565Uufa9HXTD564nZJ7utNO+tTTeduQ6SzwySWCEbVEiNlK4OTBppYW3VT9G4oavbBf
SPBuEg2iRrUyrwT08OLuECQ378qN9836ie6vfQVP0iX7VKWwQ1tscDak3IcNKOYWxFoJaGV3NJjs
GJc5mI9T9fQZn9JirCbbqwqzTSy1SINa2pABwyfSLdL/J4pFHhD+VIIG2iw0JotOAJ68KwXYCMrz
tcSiKSbwsI8sN/4p4ED30TPt0Si3/S2G021v9H54ivpkUyUab8+tGvSmY7dh9lPQZTx4uJuMaUx9
4iHLU9LL5xMQ0Dc6K2rGI5a+Y4HLws1AphIFtUNWC7YZHGnU3Fso+7lE2ToKxXrtkpO0ZyuNuVbX
SIQVYRc6N0gpNJVyiJ7CwmZ3E+My7hBH8LVf917gOWu8lwxpSATUKDAgcgh131hoTUkDWk8QbdZm
pxBcJ+qPh1YdQ+8/S1a1rKIEfk1LvdzuJL6nfPl4nUhOWpKWgT76BftzyW3cb8ybkfUbnRwBUekP
hqMq3/AdW0baMRHptOc1dA5cVEtOosFKKe+Zcbal+alaAqqEdZOoROyaI3Q2vrznhnOg/erPtXku
XkoKZelOFf1mG3zPethLQ+jOOT0VedBqfyK98vaAV98uQvXkRIRKPSlWRlmdc2WSqmo8ePM7TMUt
65qCmfFiWuRkIylQf3NAG15XeIbt/UhXm4hX6FLuW1Phuq9yVawK4YYfDDI9BDdOon7hK1c5vG/h
7Hs+8Bdm4Ta5cUPohnZW3reacsX2p6ric0s5WjHLRooY7fPBRpGELONTtzAx9QafppodUpQ6Do8s
LhLmEG5ZcpP4yiTNXoLdenDPjKS8LGsBRVGFCULi037nDV1MpLhMiPT0ViC/V6XduSerk5OyDkuF
IMXyrZ+8Lw7nL6V8FLWJZHEBWIBD9yUSshrxbA2GQr2hZaaMowhqkKFtQMlVgC9qv/OPqZ8siL6o
hGexKDsL0s1oTmtxZ7cyrUe8s1/YKoEV1IbarvZymTlFXbV0WxTrHgibZqUrHlLfFft0V32auagZ
nBNQ4R1M1JDlUpwQ1xYZlN0Ql/dR4sAPDQ+p/PYesVSBGelDcgwlle1UKt9/5FVR2nZAJfhP6U2Q
Jt2cr37w4TYIly5JYkceYpZRBppxPGWrfOnH+4/DzolooRWhpzCgh75hCNAu8SZ6+/HIOGga3msE
K9JQd47EfOdx8GQg4uMb7G8Mz3LadSohxuNCqcKBmV3Mlox2JHkHBPcke6608y276TrUvOiV+wUx
rQ4SE9NRHB2gdLm0xVZrnEWGoIvr6uCwYvjoV8CnHPcTMmavlQuLw2cOvY4gPsAkeDe28QOf8W9y
i+gU22gCZwtAW7RmVpxDQCrIvTAcVHFz4jFGSAaPK9Q6sGQW5/9v9aRuZnUpCaWVjXQY9B1g7UXk
zMN1lyq/oG6jSAqjTG6L1rA/8kgJt7UVEQ4ILqNuGKc60k9gKQX55B0WVUz+6n6brc8IeTwqbaGc
08V0PvGrmdcp1D9y9DhPXRJgTX11qLwanx5Bdlh6lpfBXlfqO/n9mDJGM07j9oe06d8MrzhiYlwH
oDS5pM5NyBwzSUwoEAj/vxQoGGhHNso/vuc4MXF0b3KlJXRui1eFebNpUDrKFb8A1ayHPiHbjAxE
jSDT7jFIuxllxGuw3B5mKWjzX4G8NydDu2sx2cQChAQ4fQ8q6XVQrp8r3kNBKEI7WrARFTBqZvJH
u41BLX4rdscbtQD2ocvoicPU16Od6nU5xJ2EGeN6upd8CuTvddq1AVBCpi+ptiRALc39A0JqYEH/
6o2V6Xvfo3bRmMDQ7pEtw0B33WL6NOc1zp3Yoxtrcjfi3LCaNrzJ/V2nJCp/VCL1uOLEzMbYJYU2
2vNMyt8BX6aGeTocEAy4ZX722BGJtRAYYCxeBidi2g7+J4NzuFceZjrbHR95ENnzJb93MfVRsDAe
I2LO99Ej/uqFAAY5wfKEOEuvKlWBCvLPapG90Yhu7LTDOFx3Yfn+EJuDIngRK7jXcvXCVuB/CuOr
PgKDR6SpnIritk0j+buqSHwXQBpZLYBHovKSzGHKaP2EYP3vWTwAMzoeTn/4hdLgLbvoEPVdBDyB
xbp1CJPnQH+fyjwkfwK/lkZXGBnmbXFc8U4HgKoXO2ZDoPM8KeUlYHGWn6vqd81/D+ViyhN+8fdl
sobK90kD8X+W8PT0fT2RuIQXGwkH7pLyMityCWBpexzrWEGk+aGDMvsdJlRAEnPK2TTsUXiN2/ot
0Hqge43I++jfMAchYjtdNdu5i6UkjWy/4PPPTTLqt2y6ABgjj4XYxutpl2FYXFgiXmh2HGxppoaz
8NKhX2ALCl5n4cgl6FomLcqrjoYZ7aLa2FOqitvKp5iRA7ewH4CscrZcn7NgffjpIaQ6GovyrLpa
WxOvWoXI75geX7sJhkoE7x+tYMRYgoKbkhptqxdzHjatU+b3Iz/3ZXcRx6gfhmm+RZN7VAGjhGr8
rYtwUSgOgGAKyAh9DQ7oRUfoNkxzSNLZv1lk9f0NEIscFiPVknD4zkknjqkkQlJ/rGcsnn5ZFhl0
Z1JFB4Xuj36Br6voU3+pVuLi5zplbslc3NVT6AM6VAIGiKSHYpwP9okYevaLO1TLB/r0HCCrS7G3
ov7DY7q67mvXGpsTo8jnZlbnV5YhpZ9miuFfytIUpchvmAbGwtfszxcxqgesXGM2CkqZMUicHe6b
fnwaCCoxMJC3FkpyNSatC4AIcTrvecFEPFG4Ayi69I7WVY8SUdDFKKZPZaDU3Zea4reohNhEcMAo
Q5Q96fZuOThiGnIpTCB6a+V408AS7sdh9EhqLd1pcozOsJsDGDA7z1CfJe4p5oKRdTu4FOKwhqDc
fTeAKatMILQi1Yi5gIVXVZqdsZXhKgxHNVExpSKIBJH7EZfdVgejEQtxK1EulfokwwZ76XnjzHbq
WWtMzQF8Y8W9uzUHkm5ODDDDT8hLTc9W+sgSJOaJDQqUuoCFiqZJMBYOnrruU7RIweQabU3bVEkK
rK7AuCCPtgZ9V/smUnbAldcESKgLRzi6rrRihus0mqYufoCSoLQ4j7GRJrcgZLdBv7J+5LqpUrFf
evqhOd/ilC4WAQ34F97ymaEUB7YvICl2H0UpZbB9KlUzQbVVkZzEpqJ1QJVgwisFOKpf9iQGxZsq
qlykuzHlpPCcQ3RfOZ4V/ydO95Vam/6dOlrClrQvsbWSf+NQyITn/STJwnEiBf6Cf092xwOYmgFt
8uQJIfUVyvvCDsB4fRrdJX5oCYrQY8JSVL0kjQseBOmuhp+pdqYgF/Ysz90xY63A0BPpmpWrMUw+
pQNuikZ3DEbevT65FDMG2YR2enPhZzVqSDRX8EInNwe7mlRmvNsVIRVNBGXcelJ4OMCOvwXaWRLi
xrNw9K6GyuG9HuxfaYtqhCk8pdEmPtuiaa7wGv2RmDsUaHVqzRX1lmtgzBezhFsomVtmFSM1e9K6
Q9V/cuF059rG6LznW0Muad7/OHS4k+6SBb2/QQ8m1qD0b09tTY1/adzvyJfnptIM33yHpX22KI+j
mGB9yIAsUY3aTrO09r9JMX/IjKjKBIipoArnKQ6/WOmPWdSHOwWI7L8mXigwwflx5rz7qTl4r+JZ
AFZNd9OfaD1k6Akd1n3pNrSZ8uEtWkWvxA+eEVWNV4e1+n7SDVs1K8Kbrkw19Z0BkVh41NZOJm0c
jfyegt6QLwvzuxZ36aMwOf4sYvjy+iPQW/H9b+Int271dzcn6K68KP7JjHtLVVRQ/miFaIXp4JDD
QIBrTviqen2K2X4hMF3nGggAjpasHIh6q3hqjDKTa9MPmZNg2C2W4aMf7YsdxbxB855H4EFQbE4/
EYcd0vQE4TR9JVb74X+HpjXq95RmfAEaa/XWHsWk1f+Ej8iD4N3+gd55wdQLy9HKcsmiDUBXZlmH
zcBvxasF4/RDl+zMA/HDfc/UqNvkLvRaYlbH1Q1CZfKaWlhwbUue6Be3R0pcbXE17AZf4lvpGJy4
pYZAeIrjK+kvFKHObRDT5EimVCwakQ3euCvKlIpJoFXDwexhm9siaCqkfM19XkO5WbiRur2RScnS
FoO9692vvJCiExtPyGmv2dohhLLOagRZ4G9KFY2Ynu2QUgb2IPEczk6ugb/G+IMaGBYVv8c1DQ0U
A8IbRzZNgPd0mKSXQ7nLYfnvg2s9OVL0IeeZfbcKtr0GGLCGjAg6d9UmpdFboJ2vZm7Mx/uliYyT
at8G5cClM1JGtgHeYVdG+NDeVuIazjCxYYRTXQKRCUwxZUxkiKmwZKZoI8HaO7tyP3+vZVQ5nLjY
Whk/4VXKIVXmzU0PLAw6m/5m1k9A8Il1L/om0saNrI3l7Nd1tQoQtHUAs+fPn41S0y04qShH/0Zi
THSA7AL0chZ7VeCDO3Vt0GY6/allVOVAd96SMgjll9PJupeeke11EzpXS2Cl7hGAYJkThotn9WGG
jb5OIOFKo+Hqp46HYxuniNDVPWF9zQ3j01cH5OsexOUylv1UgiFNviI1mqO0DRGehyL+cVcv7LGR
NWwhwyPlQRqD4A5W5RwrEaeQzdhhxfNGvy7osEw8ReINpPaCfZpqvTTgQanD7U4S7LJ0Q3G0uPkb
XThIEm8/P/UR1dSQiHGnrq19f/93AnQdd9gbFCacAITPIkHl5l8UrPvBDlg43ayZh2f7B99HQerF
wThg7r8ubHHogc4a557wi6oGP6DJzfKxOpiqqjNeVy9veCKERi0oeDvjRDutsa+AIQcjXu1AmgWv
YrZwUOibqnGbslvBeGxoI+9VVdHRoeKMhLPw7pDgOafiT/0y5lZE13VUQvKPNRWTLVFHQ2KKFweL
BeilSYsfGslmeQXFz9efVmprRf/fhjSD8pO2Btxcc/UqfeUP3w/EBiQxurLifhCr3dKv7ufb+i7s
3XnM8NMYzLsoNZWPHT9Kq35RwbbvH7kZWcaZVpfAVlaAsGpH7E7FHmO0QjOwOjSBlHl/Ap4rDMdd
uZeWQooQYHGszWHqbET+9cx7bqA3YqwfM6AcXQu3BgmpFfJgUaSwEW0+WHL19zx0JQS41VoIttOD
dLmzuOeGEpYHjBgVvZ6fJQ5cFas9TyOZtTG87lyNmz3FTXCH/FBJJKZYrc5nBXi1KkzmTG+/rlga
oY0lyKpq+9kzPCy8wAMX4//l4i2iaozNybPQj6AWFRVEb1e7lfwpzH4PhkSgxU0qHi+FmszyMjXb
Sah26PcD+SpjaBItDXEaeeKX0G/jw0VajLGKyoLe7G/GP7gB46mr1lZF1Gnve5/T+ND1aCNuebV1
WTtR1N5fepqN9/CzpYftX5gTebFZRCrzMRxk+n4nHPlr1gFBVECXLWoMaIdkIK7nw2kTy9VCNvy3
J0cOSZ32vHo61EgRWdqh2qLMVV5QadwIeCCkmCfBefIqMEKJq71Te/W6vNco97A/YnVnPF/pKGUm
eis/Aiaro4ML0Gqs/4kK+4sYDYrsdc4WHwcYC6XKyN0O6HxFhlPBpJjANPpBepA/l0EByma5essb
7mbbVniIgc4DGbhm3BATehiJQaexUSOidwwv54XDLOdvilSmy1BlHvIgf87j6Sc1rJ/TciNOt9Uw
W0tOUdi0Vk67Wuc7fMV5Qo2k0DVvimTaOS3ioiP+K8wKDJJhfMnTEnY3fV3cVtbP0uJwha3G3a1m
ogUBmF7lEMJEh1BMPXf5oJeRQKbFQSsaXk+YhO12owYja+X/TABLyJJf+D/uqKZ95l228X4SkHJW
f6erF/aG51ManRjNfHCmfqFAqsXF6MRK7EEvNJvRNIBZqznbsryUcMcXi5nn7ySSpvIMiHXJK4gW
PeC997iH/G4Y1qrYl5DQQCpIb8cGkk2v9ew1US762LAQz4CuVVEjLSIdVg8IIgox699WQWFdaBZp
g+eAMHtlIAtnSTECPOMeEJNep32foCOYxXRL8ELh3baxEqMoplLCFSTUGSwJD28uWFAdRNt8p8t9
FJdButHxfAHJK/vEKW5eqKD8q5yKAhZU4n9qtvcO6EkI/gIl+95RdCBdg+83QPQW0dvHm6MUORtb
dfhG9lieYieg0EUnYmPFX3JnAxeYPXstSC11bbmmVobHY0D4tcqSbCM86AterWpUzTu5Voiaqqn2
3YarOEsYTHgEfbBdBPvNcOz5RpikkqURFo6e6sILy9Atit2ZQP9nNqu4YgRHwtU/8ycp6ovMgrjL
y42lMWLgcSWImLF4asuLgaCNRY5fQH38WP8A8mVvXq2zP5TcA9w0f64R3IAaqFX+ZYDGEWnbzvE3
YXerQXnaNHOwDg0OPSpcN2Pj0HoZZPKCn18J4M89uYddhH761F0S+84SMcryYQZY0qvHbw9DiAq8
TUXIrufGv3DEgf/fnaP0sAadb9GGQa5DUKcXSujYPxQPGNo51wH0AA4TcF4aWBJQnrGbeN0fejru
KtxzgqWB1WPNdvfXE3dFTpxNE+dLqpXMy76Dk3yiohq7p2pX6oxTo8m0WsTgoml1ZgtyiGnrihbf
bqzEZg6pSJuUqWv1jYSpUHDw4NqcQFAWKc1O59UE6UHduYD/jkhf/5u3jTd5HEfGjtK2z84qqYWS
dPor5WaXy8Gb1oC/wPck4lMWWlZ53oaRTcqy9xUa/9JMbKEKmwZrNHASvVM6tmYRLVdWkqEC6ArU
5IOXIjqxtZm7QPKcMYpmm5BxCD7OUunMrkj9wiOWV1Gz1MjmDlCGAxIxT7fo604AM3waHTb1ol/w
uEPi9As6yj+9UmB8IrvlGpfxQm0TxKkTQIhdF+rNImtRPHS5PRWAY+N2BozRz427xepTk+kQ/7ja
fq3TR/vbeeo+z9NFzCW0T50xL+AmAPL4FjySdIAq/eRYv5Nt9c82f+eCvo2diTq8bKAnGOm6z8Xu
p8OeCOCmxJvLtj8Rg9qlLLBETFmvbF8EksxuloDW3+0Ugf1STJRbC/EctlDfi8Zu4DBXQDOK9Pli
at2jb3YPfOZNGWR0pLOBvoSP6GsfyLgTbFzmMFGUEfAx2u+wnN8nc8S4uMNas7AYRqBSiKjofqUv
qpBNSzgG43O8/9K8nf4VdBUUTJRPqWYQSbqIQcMMXw89iliboGYvrtOFykm/RMU8CGDp+jUhBUPy
o3IN1h7BWBsYUtWvLYqqitObF9estgppn3u+jbj40IlveeyFYPX/Xa1MF9YwuH4b7KDMm0GF1Dqn
/ZflFIyMUBrcQBAoo7gjNMgBAhatdGwCiDnqWmL2CODHN0TAHiUa0t2OUKRLAJ9RiBCC2bb814A6
0lQHe/JrN8ojGQ95Se6aMXyrBxUj0yV0MrNpK0SCeeeoWVQBXpx6shfy7MmC4iheqg2uB758MAdF
hkEXLBlmfPxiSdOa/76WbLhu/cpciSXzjzBbus1S7UfOUZdZeWqs/y0jja0QcgMEDvdxZfNeB27o
d7BKKBo/0/ORNVmq+w+iwRaJTIO5sgfL7UlhU2NWouPgxE8kiG1xpsM5ybnRLnw7H4N3R5sEXPL7
9aYPT/Eiqt9UAaupm28/68SkDIQIvXuggHR7aOKiwG+hfsg0RpPrWdNh+RZ1i5M6m/s5uyaS8ZLk
ewi28KYsE7o6qHJ3P6wwXqvNok5LhFwPE9EBwknDizQSwB2bETE+vvy4577oIe1njEF0h0CGPP8W
ZFkikeWlbarsHTbTqOIzVsru9Kx8wizyWJGUGLqI4QvGf8WCDev6lLLH/60cWgritmUT6rsaMEaT
/bKowCj30F5JOh8wPjRim4Tok7dk/8c2ZHSOris/gshudu3q8iy8MPLCfvlcmyBLJujTOkmDF1Cg
gzifL47hxCZCqG9AtXY4GXFiQ4zyEoaKQDjmjvDjtvoFStL6MsHDwATZpmyx3fWM1UshNvP/ajHq
TKNGSywvhWtHQqwlUcrUxEAcDvQ6WXtfEUNEMNSDt0O04/QvqoHsVI9X+vIaR5EvfMTSw8zStXi0
FUJyceiBJ2/dgRYVS7L3+d96n+JjIyLJA6vl/CY36cW6pgZwX0pe+t27B7GqeUcO9/JJgVczxZ2E
nAqTOUDu3TCi5QH/wCw+z/6fHad45IkKs0NZ89fqHcPgv9d8e/p78PS7Iwa1eDQ1RQsdA0QRsaYe
wL71bc9SsokSihqZM7vcKRkqIRGmwY3UXgVl8GC/kStK6dltRqqriRr5QOMZUhfBGTud6woUaPX4
IcnqI6ZnqblP4GKN+tiUyY6B3r1ijxMXw38XFjnysqZmnTAmq75xEX7GiEQbeb98ZRVZjwGHHEDu
oBmztKyxWkbweVcN6AK56gLU0msvy5nEL1YsMehJQOs33lvHIc1bmY6i6t5AhA7A+X6Ha936jH1F
XNUHyJdfAzsjxdacPxLsFLggLFFF0Vm0kViY6++Mf13PAfjlgseDcoOvqgAKX/BOkH1vjsY9pdmZ
SaWQgRRNUwWtx7h2GEiX7+Bnr45Rpzres0ua2vBLJ2o41h34+ULknzssh/94HZTQ3ZGcKyctZN/K
NieFWTuMgT6C/8LHw3IDTmRODI7bgNbdxadFUXbwCaldtS/8umr6ao4vl4MPOt7pY40Qe0mHEMUs
nQXTBZsKJNtFbv1fpJ6z72nJbV38GLGZ7tWM1EFQd/3EZMTcVfvL0Dy2EggWRNRPJkgRGgWbcrXb
fSqBCKx5eIUJSDQnMg7PpV9qOEpV94YwbUYoCqqqOtZldCgSkUw8yL2ep3bXc3YJcZLKgpACt4CY
3qMt5xwt0WhU5Bpg5TRcHbIsp2XJAOwnKuJOGskIhUxRiTq98FudYrPwFoxFBz+YOv6rnpIZ11Aw
j9sYyZktjOVpQBd+JFdyOWe5qG2ADBNG6ei2+b/TNIGej6dLcmrGofiG2KbzmHoOo6IzegGcNQ7e
Bx3hv0n043d9R6v7WemZNpmMZGFl6irBwg4szOZg8H46BEVQtvHpVoDpDURBBZ7CD4EPkqEl/6gP
qdsX4k0sSjHfiA1qarzhfYLSwZ4C/ITFgYHTDkKmqzHxkeWdr8t1keEqQiDpm9WRxE/jM65DJlaD
LxTYT7AA0nIKKnrgNn9STMHDSq+/a+RMoBdL6oIa2WbaQsnu8E3VmVlrCIMLoOu2iRohh7xrjbZa
xPdNm6k0eJRRAHgScXlGwAdidhK7NKmsobbdyhFMBckLEvb1hp7tOaZGEV/4wVCbr/+nCi1d0zxh
DHKfbhtU7lxu9cbb9WE2Ge1j21D8x0XGXDSg7Vw3gaztarbJhz3Y2Z1Ec9FCBKya/gp4EzAkmiz3
mpndqv47oNJ3p3CChgstUZmBo8CM0Kn+t/wu0A3wufaE6RDyjDNeW6wAPnZbzHpRwXiBABQfoE5p
cBTPlbUeOl3gJ1obdR2/+VSpsZgFRlvdxkEfUQ4+sx+v7v8VKvhGEW3DDXtz91zrfjWrpvvTM8N4
QJef0O9VZSF0I5cGZuMvWFw466HvZnkFKn7YCfZWr2y+A+aHV2PFmhLK1YVENrskqBcpScTO7rK2
ccyXYx5O0/4TG7SLeaVQ2jQ/7ycEqKGE86wMQRM+B5Te2WR8lQeZ0NlLNHduC1UhlPB8S2Z6tjC/
6x6Nwx+Q9Xde+Wc7ZwxABaW8B+hwh1u623B8iypE/ra4i5zUsAC9a3pA6lCbbtUyLqtlGdpKpVg2
wM9lu0jc+vTMN2Wh0OT4PSvkyfLFCWiNyuWLL1KB89ojbY+0uUEhiUNNb9YSs9qYnhU5rLERAwpl
LgHFZjnG8JoI1rB6KQsR+RmJRkzkdsX2Mgo9lkFVRDf6zH7B5ucwyUrck0VFCEDPVDyT8B4YCTDa
W0JpOGcNRFBsIbb2VeekLJeOFpfvWKpnXF4y1tzYWDL/JsVyLI8VLsPAFKEfapU2aeGR9+wcrg15
MOyY1eu8EF6w0g+sdVi2ZThN7K7qErOOQ8X2mYP6lHafkDMBByxErWc5w0xTCvh6Ss5vqOqM89hZ
BlOKNKsunKZBXd2uTvh/E15fWaiyzrAjAr8xU8X73UB1YMWDx6FGMti7SOb+IkNrryL8FPo7ViG/
Uf7KKUu83lf1weLnVsRSznvzySHGAGX1m46dYjdyUocYd1fwdYBvJrBMyuCcWkBwJdcyxIhGIuSy
1bWjwUbgXwk1Kw7oNjPBew13I3ZJqherikz31SgpiB+6GN2AwBMvsxFUDVEo/a37hmYvkGK39Ww7
eDG+n/guF2KSX0Z/4Oa28NDju8oC6mb5/rrFdYrXpuyU18PMBhmVgOyFYmJ0Uy0h3JvwhPmboUv6
dO8H6kGTZZrg77qZ+h32HhjFrsE9tZH4R17RO9S/4RkpaBC5rVx87XxW1+xEbb95p9ywUxma018/
GHedgcm1Ym6FbJHe0v055N2sBezR0Ck1sGT/uUQuGYzmPhE2VKU24bWnDT+ALTiGruQFmg+8E/uL
SONb0yIAcDtqYHuFUk6NCvFKZYKnnUod+j5VTPOlD7WElOWklT+LH9I5XaSJKMsopSzKf4mUMMjg
85iu2RwOIsAZ53miztXnWXsYpIBsYKgoyFiOYO6MIFY2A1RJ9e0DcrX2i9e29YIdUpsn0Kh6V/Jo
LZ0pDjci7nheGg5oTDIiF076+1AgVdERYEPXiEe6eJcF3XUM7ObLT+sTDKzugX4fsT9XJOPRFQLE
VQJSqstLww7EiSKp77LGbGS4Mi/kDCxi00QSolvFASg/8/OU+kJPH44O6wEaptc+ZiKA+DcphKAL
sT/3nzoaQ7fz+qticah8mXfJ9Z3RHxoEFFWbabriSyl0Xd+u5MmO6Id+B06kTRSnecFKsBGY5BdM
eUYZGCZnRlmPqCR1+hcoaqkOOwnmfgcCl8EG9Gz8Q15UfMgYbkNil/2rMO6xw0YsIDlN0mE5vmGo
pBSEtUUER5a0DbnhKEMIykzjxFQcBlv8S83J+G2Veez0/1Mp0GK+xhQCPE8/Jqi/t6JwBpqwgHAL
oC1b6BzCiptp6egaU+fze0iVAXY2s5AheJ5+RAaVFJ6WY4bk8cg8PUPghv8uA6srcFUJj5dVGabg
Wh+Y7EudwPQraCWUvMM1mjoZYQ9xXWZto2NLZNiyoyiffMqjxD2AUMt3pVtG9Nerryx1A6rpxJ8E
qrkp0vaFYRN+4ys5avKGpRQ9rcWbTJn9RVNL5KstJhGzUELerfj12DiwsBjaAVCk2abK6K9ANwYg
o6T7yJ7ZuRKMZ1wVgMXJdvnwuc4V8NMk5EKjlI/ZwKPCxPLLIt6HjRRSXb3SAnBXfE0AWXV2qKPL
NgFZG+AkV5aQzUmKguMHIFbU3MCCFI6xnPLy6/PGiuB3e/8WPMArl5Bur8GtcIIgXTYQ3nINZG3R
CuvxtbrY2/jnDdTJ1apRAfp88c3oKtyrCN9ahI7t0flK2sS7ngJxex/5TkbwLZ9tTAX3QV9BebpC
3jf79JI4tWiy6cplGi2oNMmNEPeUxVCUFbymPINJs3U64yy7ZdChb9kbHPwRhGLzurAOahkkMBMf
T0xHlgPcapv6aQdrecCkSLbopQdjT8pkS491Gyl+2kEC5ZE8pLZIFFIr/AnDYhMa43XhsP9rSZbT
kvv+VVTYHK3f88411wAnIMAur2CR38e73bkUO/ZsfFhF/XcW7d1zSd8a8gile4ktmf1hQkAnChpG
3w8lz0bKXn/5Lkciqwv+NQnOHDAWwoMZtI1/q/DhjGCKsObTaQbnLd7Ye0zRSircJTI5fiyW+rNA
uQ7DPEyyxzslO2y8DH88ncP3wiJMSj3/9hWGik6MIRNXcFiNmSEk4GIWtsEZ1phd7mJ9UnH3Sbqu
IKD1ey6n+mhjTJtajBYb9X+DuDudlwC5YnzthFxBC58UYdzJfkbVPtVTLnu0sXspfqJ+Xo6xrNID
HSji1Ce/hfDWLCTQeYIMS5G5k+8bY7XIETrNaM/a+/hXa5KObo84fAR2DHwIE/du7cnsZcHEkgTo
b/2mXBTv5doR6z8SLRHQtG9rUppTXoaUSt8FldvDDWghUOMPYvHRpCKFget0oyiDPt2wL/54Ap1t
BdmF8YEMaKGrbSIq2fnFwoQnffQXFABdHg6YYoOhQ4tWrU+/qSmCBbfaRzYg/Q+aujuLtlVIQ0+Q
WA5YK+2X68C42l2HV48Fw7sC/8hc5dGLz4ZcJRy6TMP4xXbbI0Oh3Y9oxhTkxAbc7W5i1+HJWXP9
i90sGwMiAn3mmrB9lxqyz58Zg64ymYDXqFeIN8KX12CFqZfWm4w+L9XRvHLQhnm5mrLXWNsaiq/p
Q2BdPzXU/Zxqd6iTOJgrihX0X9bIVX61p2rMcSuE51uQFtPGAs0SO7vMKJ+xxzCtbcBXpRzzOmmw
59f6mGNqNwGewhQz5Q1G0ZW3hLW/cOmvUA3Y81m0rArbQd9vg+R9UG2YHOz4q3GAeFD3HegM1CRb
CIruBEBQnDsiDR6lDWWh6SSr0dyY9DbDQ71fBsTcYBnhhbS9Cuw7nI8V+l3VfP/YPlxlbrDsStnJ
SbihFkqlb+y0aVi+Achj0rGopQkP3d1dXwHXPt/IInrpb+8T8D2M1x0qxat55yxQhpPvD6GLeMVE
wE2X3a90ragX2QvrQ6f1OSVYZIhlKoLZVKPkvPCO7/F0GaFJTjtDGhXNgkzeLLrY0hmf5MjcC/m5
Fcypm1UKhILnVoHFMkAmYN29sQN42FfIg9MWAUTxynscD7pJmOKSlQ6409wB4+LZcPqYYfxiHPXn
gyenHKutSy+87pDAGTx0CjPc2f9URwPJbaBS2OrutN5nPhO5tYeAegSrj6c8gml7Ta3zbZp8gWmU
hytXlGiJh18V8zS3I5vs+X4RdSkg4VXz203iKdP5i2jLHGfJqF03yinHfgNfNItB3NRJ2gWVYjiq
7gr5bcdY3fOhsdaElup7H4xjxI7emJ/roaWlVb4VfxE0tkrWfB6Ol9dnd0eVgBLyb7PkJxzMJMmm
UDykDzR+PtXTwROhQEayBnZoDSAIPkkN4ExIJ71NhF4fPqkMlc0xgvz9Keaz74k6aet+NcqHUuLC
hfPTZ0YAhSjj2NUah0OO76oqA5rhg0KWl1LwgDnEDQh0/8y9dLhO6gw2JYScQ1gicPLnaoHHfRu1
3E92UgHtLUzbvOhIgb3UJiyGidKYoY1iSzE0Ni6QVLW0dg3T0ASr2HoV8rhX0zrU67Y6MRtA5urm
ICJxEGlZl5j83zC9jfMaoUZJ+lY6KxXCdB3uA9SFQ5vdaV2n6SV0hWKjpplz8v4erV6kepZTB1jD
xiVPenkN4azDUmfqm959duFlyz267OR4py+h/TwMtrNuvPkRoJapYUPKWVQw3jAS15EK6z05O8w7
Clmp0BB1lAmYfzVDunbBPj0Qc16N0rFi5jSRme4vj2bT55+KviTQ9u0k4wOem+s2i3vwUw3w+6hI
x9qXHxh+fBY4jFJE2harzMPG/Yt4YM1MuJ+sIEofZBIh7KHgDnmEnY3wuZ2RWd98f6PGPvVcN0Zx
rmJ6r8waX1nZ8l+mAFncvTUlbDKA7MzCIyVRJPcZTR7wYWXKObgGHqPnanAeH07XxGuXrSAyIrab
MSknESiF/AhNX4d0hfNMNCLqWPe98JJrPZA4n8d+mwPEg1TIufei746CV3WbTWp5NttZJDqa0plG
VxUuNNH1WNy817cPo6+ZrX56DaPboDDoLfVRgQdTBQQ5vQoktoy07vUXF8AKLnOUokqlHmnhB2gj
VgP6LBWGLLvTsV9mfzLRPVgpP7u8mVE/xqv2Om5/IL2z5pSMRJCZZg9Q1RRFN1sDkZw6m9hww7xz
l/P4DDkiMzrnf3JXCEwJnIaZIrNCvJpvE7qf/FoIUtrWek1pX/8taVK92Y7FTzVA7HFipzED86Y+
P1gCAbM9OecXYt2040TLugMvSAVTtyPOJChlIWRnxA3nSc+GXNS7NDA/QhlfZtkzfFbMRgRlH0ZY
COtd3mWh+BrXBYHAFSsAEsdLXgVz7ib2k9ZcBF6/GWwUHkNB32gd0+iA8sVlnXPehlqOiGHmupyh
99zRFN2ntkc86T88JylOcoGLqr+tKtU4m9ywSUnhOwSbTJtrjmltMjETLFwDRdLSIwVmFnwLXpPU
c86HApphWdODKJeqRnw2PN2HZ3xKL4VC5AhumWU0BG6PHebXFC4ev6pe8zMMMKIU9ix1DBy3D5id
/3MXeaDGBgo1ZSn2Z8itDo006kp51ova02pCHoU1R3vWKF5V2qbi2hiTRqh3+y4jRFsxiiSfvl7V
SjG54BvVb1RCRG2iOANMnNhoq9PJFcFUKIG/b/FRwsYyheX2vTvTkZ5Fc/qbXFqn1bBeQ0+qsih1
u/ASNz5LvnROKJFH/R4vqG0z8QhCavdoVbyahteRIepKe8Xcddt7nRlRxUtlImGsKVunt+HrzoOY
6qV3vY3sWvKl2eWqRdy8hApvBrD+x2T6OzTwikNgBn4b1Dc4gzfPGfm1hrges4qsfoj1hMojWyFm
SKZi22SYLEiHqo72Q08VhvpBAviMpHCGX3irWF2fRDTDZgIEE1nXorvzMZBO0smFvhpxV9t00jlo
FA2D2Ntghstnf0tgWkER+yXfRRauvC3zMsJ0X/6i4igotX/+f/VgbLlRTmZB15eh4X59z8QeGbSU
iJ/cmRX1O4pP0PyXwnexr+tVi9Pr5IZMwzGR21xXn1D5RgIrrCNLgWzuDZG2sg4lqLBV7lThxj+o
P4q9KF/YGw1Y/kfyy7E2ueHymUjzAZ3GV8iMlrnGhZtCxWRuB5O/GT5ZajJK1M9kb8BD4T5RorQq
vmHDIGIOTadjDN2NzbLzac1y/sQAiJyrZGI8GXES/VYuJJYh5SQS9sCGJXQuxrFsx6xH5tq2+CI5
BshC5Jn3vKp/B22GJtbWbpt71SN1suNlS9I3morKBj9XczymveLdqyEi3NDXlWUXupRF7pQQUe85
QgxSxIlmgrIYqnTtWnPAbvI5AICknU7+fOUZ0lkVtonJmIGQzDbYhyVUCH+0iowcBu6X0ljrlF23
dz7kd+HwV0RSx/M7JtKzZIbAegHyTfVLqRbEGyFdzr1mjUhFsXbd9PVMmddFMWPTVWyOYv0SnIqz
zoHrvDVa8NUburgZuv+EzGvamBD4Ne+NBqrgwL/qyIZSiv8SfLcsh9WqX49mWj/Blr3wUm++tleh
OfSyG1Ya4XwbKu3xwpFwDLKKmOlsJlndV1L1uDu7Uu3KNdzGK1ETK3P2of85jj+mWpbO9PzASZiI
9wNm7Lus2dlf44qwcp+wuMCHZcBg7tA1lVb7YqmdKPsOcwNZsk5LOCGbkROgVURGgr9a/bNvCqgP
LoM4oFoUAy/eMA0G4BTYCoue53gvYdLh1Efi5UtEevDvipc7U9KYGTT04nYvZpeyL5C7oXFs7RqC
nG63R6oWI2JLDu5jYYQU5ePJs23EXKRY8B76975NVTKXKJQQPVYVwdTxJswGRtRx57mxAgrdv6SC
e8tD7JIJywNoci34BCqsJcp89xtfMFnw4xxj+WcdaLOxgsjN890vLMooq5zsOZHNL3ZWmbupYQ9q
hBdPFK2w8cm3pXMUBay0c5YCITMrkB2qGlPv2aifeoWKN3WhXc2UKzWhQw658phf64TrWrhrhdTr
5NfJTKbwMpMDdt77y37gKRNdIm+hkFgpxgk3og45ar49lbK2wAp2d40g8A7gmIJjQm7GrBdBRLAx
kjuepFL9x0x2uDxn/20vQ0Yees0zEDFBqK/UUORG+lMdV3957kX3HavclTGk2XmKxFaG6LkL5kIC
+JC9YbOl0X2R+2gs23jxkRAxmWJ+p+lagh5UUm3N6xZ2jxsCA45Wf29w3IiZ8EJpmb8a0xU7mGxd
CWuXaok4WYzIe3bZmwKh67z9YAGHEpNZJWi++xDB87n0ifcmWN/AP7AmG60uVmz1CKCjhBBUAzHU
m2TeLWx4ZtjztbFB5VjMFayNG5RHuCuXfRauiLpUh+77jLXD5wzm+aKEGuHievvrgngzeh0nj080
DctVnxqWg9wY1ogxkva0dvYLtFRwlMqhnPSjHul9vlL1mUDyu1roh/Pg+Ju+Mufyj166jBqTpLZl
97kfSnpFfzB4I69EVgpJ7OW7NMMcbOL9ak0IWdWbDPnrgkqTRf6bUMmqgEBBbimpUi7WE2b/pEml
cj3JrTezk9QyxANp1bM8DyVUEeO9ehvzErt8McT5ysWCjrNTjrcolOHgkiJBooljh7yD62uKNV3H
oXurHV2g2kPUiu+qLmHEpcWlEr0cA5ibl2+e5DlnyAKZzQg6+VNMKHldzMgen4u9DRgRueD83A1B
ZO00pXof4B7yc2GDtRH3E5fhSargrO+N0Y7bZurs+jxeM0/waJFRjaHuGqGM+dhszD5Dqp4PWycE
o6EAp6Vf1F7jFvamG/gOyIFJbqkjqh/kNBchthxiYaBpO4w40AADiqdg/1KPJ/jAgteKlOniYX20
bHsEG32qPkemQEHGBEoEkT3BmG7X51hqiE/21yCJ1VtuXB5JeCh6A8YK/bX7cdWIY718tOUm4jAg
Mk0dXTpfLZSGMq5QfHqPomP2yNJHywVVXzMQtfRnMbAjlNsTk9ZGYlXz8tKzeasGo0ighH1jjA2w
72PbQRSKVJFeXHLfQjjPjiyAEU+O9a1EFOCukbo7tjsT8kM4AkP4lOXqqzO+4qCa/Xs1nYO5W6YU
vjYB5Fz0x+aIB/gQwANO2OokyltEvRiWIZmx+mkQ1DBPI7baWhfRWcioMrQQWpa/sAzg3tQ5Y4T2
1XMO4g46h4UHcwMyR+QidjE9EcXDvb6RPqX9OAZc68gr6ovhIFdDz9ZDd5XXXB/Z4tzPIUKZ2o4v
54ZbdwbyVfz+UkLx/0H1i2etjxS8fj2hEHsI/GvivyaTYj/+nbGG+BOjAR9NFz1s6B7RNM0Tsrg8
A5jZUuoHE3pAOC+VBEv2b/o7yWMEObpsM2/aXwrop2EBzWIrgYRbdqWKdriMLLRjKTK8FM6OrGCg
PGEh7vcWbDI3Y39of6xGoz9CZWX0ILnS9nspryksUQ8VojujuAYJi88C0Ul7JkrG5iiwVhBaIpG+
Ozu5zjngp6rqkintvkUlinsMzBD7TsnBl9iHX8Z825LgZj7BZ94atkquKjvuhEYdbZ28so98mpoP
vzSF69xRZSCR6bu69J9SkQuKl0J8QrvGx8m+Ce95dQRc6mfUK2zi7VJMdAibgUBRcXnCoUPQX5no
Cs5Dp52K9oWI85yvAWf4Z6tTUAflZQ6cW3UAceEWBmS4iTZmFdpq9uzwDQxXhucR5dHi1Ls3jeRO
oRpb3TOiLLuNbilKy4tNPymKpsKhC/w2IUuw/NJHdt4pLfp5fsxZ7g1gVZHslxOgHiNmMwwvf+e3
1jOlW2b3w3I6nwIxpGhZQmY25IVLBzUZGaDJy6WJ+zmRMCpDAzBDM34LK2aXH7TtgYi/dqG8PkUT
cR0TkySa2yK5KCxpNL64eXCq9Vo8tUZDAiI/sUHdrTrBoSU5fXx/UyKADoyrp+XFwZ5feM3gGoD3
COVlNOu3AMBzsI2fQXO+RQrkiRfs50sdIt/RguyDZFcpQLVoshAEhC24m8TEuZMjczjscaWVfzgl
byjgaoRZ0bHBy8s7bR2rcBt91byuo1CbA8bK7HRCzumD87VMgiVsypCduPCPpX+6M/eS3J/f/+nY
lcZ6j341a2MwB5e2XXaUIsue5WK96UwDJ8dFXouWWZMRhA16ct+gYEtnrrfJpbPAeO/Lpq4aSFez
GiYP5+k3xOdHO8zAr796ZlWFLoXZVz9z50LRZhGoJd9iQLWunWbLLDjGVvmtTYQiD8/UR0QYA897
tRXUzf27u1P09wG+W6mYzqQ3+igLBCH+6s0KH8zMo2FjsTgKp2KUg35GFnLe8+U7DAocQdOHwI4Y
V4tTQAlQiTcfSk5h0Igh7FR6F8Fg1ZnURVLN7NVqEAgdylicyUShQZ6fayHsalKgjsuc900coYLn
h+aX7lvwLEYSSE4wWwpuMu/1cOggZH9y+AdzOAUi4sETTxwONVojgkMNLFS6E0vmE2bQ/UvQS5SS
yUb9YRzh22ym4YYBV9UEYM5YvxPERcMCmiz95e75227xM5JMZzoZMTxzz1aVG6/a3iYwe+JS2tvQ
BoVEZe/h7it6KdzsjDkJ8//uUhC5IozgWtqnoLPUzhNwGKfwpUJwBZG3Z6Gxg6Q4YINfkgWIRtXF
MPvMTzfsIkEAcvmNU15ZrOjJ5Surx6stB6/vTeAC/gC0txKbUnDTT7EP0v66gLR7+phe/RoqdUye
6llxfno8q01BJl+Jt/GZyKoYwSX/ntFUCrnYNRuuSYyPwrSKSgLBxwTycno3WbRaMbWJCcQTpSSH
TBIxczQOnjd9VPKlf7h3nCaLmHpjrhC9vowY8LCdg3Bu4iQPNhOLmD8lhjyMGehkbZzdBFtRObUz
PYuS5vrnrzT8OEaKD16WXuDkj4PrGO9t+qiI8lZdSaGvUPWBGN+CP25VZMpOExaQYGMKFISaM3Hx
9U20c9AVTJYpPY9nOEtTAwNkxbqf0yWXXZ6Adzm1NmnKLTvMq20EwMALs8ouHbIuuOl3HUsoTB99
zW3oqpRLrppvgH0qyKvWAqR8n70T+gnBTKfQPdxA/qXbg1kJ30ps53gGMRV6JRu6YLKUu8zsyQKm
CIvXz518E7hCVkyZUAtSdUsHZzD3Q7BRuAjCjog963FE4UD5UiIkToZvnx6XsOpJUG0bI6z4TXNx
U4waJsJ1Dz3ha6+m7txV2GbNd4P4asaFXS2lSQ+OSgaNjwNP/3+w5k5T8uij5sw+frd08nALBYWW
GPhmme6NiGH1+lnbqy5XaTP9PiBH75A9nRXYboXUG0iqfmoibHfQhzJDwAb4ERpP67aNMfT1nMKv
1yqp89bcIDQLEUBtc0VAaGdxA+azlDIrZnHhH4q7o5uUtOvL1mvHH26xasnvacqs6aEte0tjr5Sx
8txw6EfPdnTYW92Zmx4fu7vfnwbBuN/UpS9ixhaedJF3FH90Qx1nyQQcUXICNHXotv0gk06HBD18
XlprDQwAyJ2R+NK7UVkh9gK45l2faZjrXlzUHotZzyLOOd8eL08/iTkMXeSA8VYvsMu0fQkJoao8
9V1fYZBYvdBMF9wQWrKiSbwb5ethKWGSzPSk9LF2w9NmjTCNUggZ6Xap0gMuXIBVgChYHJT1tLH5
NTJRZ7h5ZQL1H4VZtgy7fJSqiKv9TFM3hqTPjAUjAMCkwh7qQqrHRPjyHBfIHMPFjV5ZEVezmdz+
ITFHJolJ/ryUchgC4M5MR+3dilt+2Hlov/1eT4Jb0lfJGUCrKPTkkcCi0o7Qx/myLCPeyxUZSc0a
Dtgkv3Nb9RooG76XwjIU9wk1IiS1o9r/O9ST+urQmqE+ZMwSWrScsAObAt4pxpFdYZxYcFm01Ud3
ouwpP3q4Zq86WUvNPh27zUShmLxVqz27v6u7jtTEtfWhiuPSQoOziIomQqZVVsHLs2K232dKAqCa
xS1bwRiCb/9pGnkj41tO3ZEREWgIsP5vnYsrN1/6HPJ7+P0K193lkMiutOewW0jPmee7VRRnU7UQ
GeKh6qicVupAewc/3ofp62x1D3Ml0rcv/X7ZFp2j5gbmhcrc1uMpSE3iUl4fpfb9ui9oCAcCYYvM
+GTwHc2u0Ga57u5aNT7QN4HEUekyosBoFzTORAfVfJzBYisw70Xs7SgvMmdf+zw67oSPbD/001/b
D5IvOzRYQpKP7Iahf1kEBt90sdqTtUqeKCcCs5BsqPfOvAhIjtvTHLZJDI3qPN6jrTllQyOiRpa+
zXzJl/hdbVS3yHs4ZTN+iYhhxdJhD4c6LPM+K3W48G8J1XbsMyHk+miCBBBtiqwBfuIjYd8/whSV
ea6/6/HlCiv16kNx1W1OtsPI3/NteFSWyfciwfYvrU1S7nDaGOgFAnC5kIhOUkDYa5mwzLmvXhMs
lUCrxwnMMi3oPAvWvjXsZ+SetqIMahVgd8up3RvrUlqtPnocVnXwCfH2GlKTrdiQShz0WCrDzzIw
tGs971YTGbiH0DKrfUjAneVe1Wn1ES/96vriyho4q0oREncc6nGLWTL5b9AwfIMfa8snRTL7KNuJ
Nc1LwEuLhxtlBnfczz/KUjobNq2JLWr3G6XcO5KzFg+UzlYDjVaON+bJM3B36vGaCszjy5gVSe6O
/F7KvYTHmU1TGD/+LQ+4REtSfumgBiUyJFuYmz+slamyyp8tcynLgCvfR35L1lFSl0cceRse0ldC
eBkKMggFZwXGlbP2mTofCEHgmgEQDh5xftFc6pZaMz00lQkMviTmTTE2srEDc+J2uQNoPZSARdaC
Pc6KBrF6KoaEeBPFFBrW/YBFAy5qshxvvAPHbZoRByNwYOS1BqaW7wansUwA7Kpq2XlfP2fCkifE
hWX9Rt7tVg2AsYblxjNF3g+l3Oht6wU+Dj8wgMYgciswVpTtXJPHqh5Mxd3geTofqa0bBjIJTuvu
zhsleDblQAsNZizkRso82pkFRc9vjt6UxKG9SHyo/0mVd5/8bhtUyoqQF7DjNWz7wK4pp5OBC0ll
wgrnoAw6E4aRptszTfWIcp5YqcGSODAh67bH+ZhNRPOp2tl5HNPG5jxLGE6SjxIWQvqc65HjE+nu
8N+5HWS7ICuhWWHxQSweOVckrtzb7lE+6CYGBPgZNOHl6bWxxvjGtDQyb+DBIx2ckI05rWniSg4G
GkrRJ+OAbUMZcN24h4+xYKSPhbozCy6knIPlTufHrfkiT4+k1OucSofPi8ir/tonOhdBIzgKnC0E
ZA0kAxxnD8H4ArDdD7XnmdDrSl5iNhyVQ2Q7KejDQi7gd53obqPtm6QHoKLX7puHylD+zJEG6SCF
gcLU0IryN+OUAqVdifYROzFrbS+KlLTu56g6FIwCKRHGliOkIfYTbhCQhSC57Asv27slkd1kemUF
HnJqh/D40UHqxzYSXwoIitRIRfqtewoaxA5PwcLLRocNtJTJC9D7kH9dlqDbcmjfXXEgutFJQxNe
ykQ1TYNE5c3FyOnDaGcaM27/Nbt0rtLC/jb4ziLujjACXdebE/5fxrxPAww4P216bYPp15ApXBK3
JRlxyod+9+0fcbXLo0ivG3tNCUFF3pHomdH4FPq6O/5R1Ps6vCRtyIB0kC+d3gC6/9di/WU3oQA8
QSif4bozLfRfVQU0g8wsBnh75M928MjJhjKTUZC/gMB+2TqivGJuS+HEceNyOnyEMVdFCLza1vHI
V/U3ZUPtAMT6AzL6wKJmQpa260HIIsRw2fIeZ/bgw2nHvMRHQQsbRrzGjNn1b6NQ2lJNu88uvjwK
xOY4Qg2glJFcnN3dS0GmzfwMKeKmggv0AGSbDhtmjiVXL/O4P8GLW5mmYzPqk82u1e0ipLQVdkBg
gcbpCCZntMwwGbZidz04+9pSuoEaUtX17AahI9VTsXa04NdTvUXwMeMRU1PDQe0MHIQZ/J+47GSc
gCG2TB0bzKD2YhZNpMcEerUe1CP1V0DAY+b5dNUMeut525eFtCgVV2QKCclkIdKBxw1Ms50e1MNG
RnWR226JNqeD/pbs0zETZh0c6ZHYWTfHVTEhKc4kE1zJuGo76AEYlkHFdZrDTpz1fosAmYX9XNDk
ZwmCOPTlwnQ3CDEYIBC5+W1jCgwEiWygb/4Z+XrnFrhG2U4RjDCEiT03+KM3B5tnfUKuAqBpfU7J
IEaRsOBhqagSC/qbJFwySmCw9UGKBgbhF7P5D7zlCRdK8zENa2snqyt1na7FzwLazj0xvsLEy47w
TZRQYx1VlZgtvUaTecXz3GjL0qTWbxSJB133eHHRZvjOPmQVAjXUpCD7cw92pJO2j90SelphWTmM
Cj3PVah+eK5SZlQv+ateGSvLgcjC3DAfmzJOyGz7guNKh1PEvy/JCWMxiZbdCXy/FZyv3m+8XXI7
Ucg1aEwKwpoXTinZtOBFzQpNlOSux38vpzR536cgoAZAtJB3i1nnEz2sPMLdGNpX/IwMJiiKr4Nh
b5551KPCgLML+NDc9degz55b0cz2hvm6EwTBwGDboa4nsdxav9ZTqNohHXrh3+AQ9X7OlzenInYD
+jiZI0PvuZ178LTVWwwIAwywRiCUn8U3JmqfOaM7GKPBngxBhXu13714Rad2p3rveV/Y9vm1R0Rn
pDdwn0jIIIJWjbKYvQ3xsMGVOqNoskTE+1i4EjOK0AhJCyhSaVZVY6Q82ndlhtgv6DK+JQejzS6Y
dJaK8FIP+fdhlKZ+VZX4b3jroSp+UW/zVdCSCETQnKvGkt7GsRtBQSdwgh+5JsLfF8lLJ6oXPpgL
rOLWikiosbe3fo+iMNCWuGh930ClrNv1MCsvg6n7FkObKLv4I49ipakNlexxXGOVCYmagdzvA4P7
r1U21yo/dGRgeFoPXPki5dihPvYpO8GNUVPInKTeXldvOOuowCwDRB7gQR8VRGqzNj98VZ3GsJE8
8PtEdCq2Ov/RfZF4cbrf4KbpnCNq5J6ng1BY3cM4s8UuJNqAScfNYfoAKloPAzW/ugNOmNrOX9ow
Zru9Iz+kxB4AnmBg3w2wxN6IOOr0PbJCrMW/chXX9E7JU6C9bTNOPKVKE0n+vX14DJv5DTklnTOO
0Fm0WPL955xUHV+29fH/5tmB9fgYFkdqwgNABifq9JdjSxkKtAZ+V1zA7oEIGxN0t4dvmapx39VL
J8jwnCnxihcZrWjcHLhbr6hAq1cTqNIrgWgGFOvm+znGom3mcijx+5OxENC6i+aAz1ZSmASTfuex
9BnMgxhaHrsfmE+otuQ+letChQNqDYeh20taYaOPQ/M8XNoI+ibXW9Jw5PGduqS6eQxMVk+jGjVo
ARCNEakKDnJyGQJFpvxBTZbkCeB5NUrfRsqEnaw34TijhqU+hEu7u8RXhxrK6Fbxl+z6tieytCkc
xkBUXpDbUORIgLAeG74871B1j8ng3ydm2i1v5WjCxtXce0tXKZpJ6r+qwgckiAytEJlYbAbtR6cA
ZBkQGQOCQvJ0Ah2vQBPFo4lLATJVlCeL/tBDUhcS+F5IOrCZyvrmxrnqoapDg36QGIft32hikuoD
ghoA/2vnZNcR62nSLGpmwaJCmtXgAO3D4fSKj1owcpD0+xqH9Q2kaiMU2VCTUTAw51NZFP8Qgk8l
hUkEF8+8wJgfWjyzyrGLrRoqzWu9zsUrNatX42t4hjWfWp2SXPZiJhxymcVLw5so1FhLq9vMBvRG
QN72XZsxFZ+nIjpyUkWRrEn8U3EPG7R/XD+MmdNKwhsiQ5Ujo5KAbY1Tg/mMLBuKhLOOWZTviuHe
5yoVu/V1/7lYY5oD7wmClHJPWCnFC6q/4VxioPCsns3/tC0IaGkIyx/nrGFmbeeDOR1NKdi0y0tW
r2O6vwzTlVOMpJhDJG5Z4mkXTZ2LgnEfx6opKg4HP5wcdMYCPgdkcsmEJKK79knk92Xyewlkr68F
Z/ibEKzJhDj8mAeBPFYL7JTyXNGPoDg/8kx2vl+P+7fFSv9mlBxgwsUbNQlvzHr75Ef+5VFT9ks8
/qBw+bvioDdHu2Zfo+37GJcrF+aRjHzwV0NyJTIfjat2syIIo4LTrUeE+od4//qUfHWn+PJ1lwmQ
0uLK8+QSrcduhjMFaSn9y6m726q3lPvmpMudvy1YjYJGg9e3d0U/1tWx6BHZwFqfbQp7/dX5d/8c
l6NFeWaKY6aUw16u2T3nTAOhIaZNDUZ8LHXvTTXqR4Kc3IBNk72BBCXt3szj/6OcpdVguJFCcSOF
72EWYTynv+oYLU/8NBhDABqn7XrCkq8j8BplMEgms5xaldvC2UhlWDJqonRPYX+h+uEa0JDZAjdk
fmQS2CkWdL6maDHETS7Yqydp1PwBeP1xl1e4fH8NOev9NAvEjRuIjlONHkL1JW6Me2kaz22VW57+
QA7s83pbVUkO+5OWHxW/vph4LkqqU+bezHjjFGvK93916kJipJaLNqvZrH9RKXKOi4FMgYfKKaxe
bM6OJ/2B0k5oY0T43N9nin+C3REnaVypjsWHgrdxwFSQ3Xpn0fGwAeUn19MXdDl5EANk1yqPdL9j
F5AX/im9pU3rX8RplpejyK7r4aitGFx0bkHCjlym0qocwegrjKObJecmBTJvCdMcNcFFV3/Rr7i/
pHkwL9r14RZtqec9H6EsR4MZGfL4gZ+V2KE8Teg1/8Cm71+msKedup1JEVw8tmRpyLdqWXRB3grb
FodCAP3ni2VYzBnAh3ogjudd0SHzeuP3kL8ckWsyajIi/HSluRnkYQokVmL1L5dyR0KNo3gqT6U7
+BcwcsIclPrDnm6XR7bYoACAQXsoiY9yQVzValpL1jUNFLPgbpbUcbLr/he1vbR2sbRElIaCf+fS
nuP6HYnnwIeEt4jxFxHGZP4iT+qd+buxzo1khkfd7dCPdLHUbjbzNuHm7FkpcnXMM9Zh+d1RG9Fe
ZdRPix8DgmH31I/lKREX9tsJbmtGH8k2XKDCvCrOE7/UPP8lOEHaiMlqZZzAuj00FqMr/8xU2Y75
WBdJZX8ut7aTWT1ahDB2bGPHS/80GlCBXx2uhts8ZbNKk5eKocihlLqVzwpeXNOncLnXFNq5mIsy
JxJJGYOJrvXja9gouY1/V4zmOX+Ka4poVnoNDa11bnRmgtE7VTHlVct3tqJW39jJd6QHtvcd2V3I
W39rSKyr8c0VlRVZyonGnRoC8HM+4SOCi0lOZyhdzUJoj+GjR+SbbG3SSWLvEMh6/ERhhwmjhxBy
KKi0ObqRbWMIVvl5XgU+fV8t6EKM0mxt3yyqNYYwSTXpVmugwRlqJEJmEvLpxeShSLOxfGjwPWg6
LExi8p1Bc9SF+xN7xlCA525IuyOqfghdpyjon1mBOPRVQWbrazvhWMe4oK22S2FXPmspKwNFmFWs
fusn7QJle8nPbGqlqbObKNLdpV8Yo9yEZL0my4yMO+NrwoBXjvpOPZN7m+p9MZNANgtTh0kPQuUd
d+VEit5jVnQYFiCjjS8iDNlW8UczPNmtvvs/etDEsMQ1Ta0WXaMuRZT+uvBKpThejiZIEdwZgKIF
IEvXQi7AOrDOF1jHt05uyud1H7ImOjm+8wL+Zlxjn5kVdb78oqFPOHCVrpNdCjVa++bfQof6Gdav
v75yFJ9Jv0rLC35gXBFDov7SYcgm+0wNu2eR24fTfaprTGotGKmqG4eSyRe871Fn5A8ugH4aGRpI
CgttOb+c5gFxMLPM3cBV81m6b4u+ssAnlPUTClzzf7SHhbA/uv9H99UBRgcUt5DpRipoR28fCWF6
43PSBPlvx36TEBKowAGWiMxLIfstpQ1VY/W07ssp33k6xAsdNvJADe/Dg8NGFocMKA1cYFvbKodE
nGPG23ykYG1w4iJoX+KaLOVCEO2X2CfYUINVOWyBWCqIPLENvA6duEkYn60iMDNOgb3HRaQZrbQJ
gOyu3Q9iKVKaea1S5zDqcceOJKuaYkDq7avdS3uT5EkcNMrcN5CtoIJErH7cT2c5Eci3TyN6DIbF
/H/GsIbQ4tN+xTjcVF2jfGo+OE9ui0VOYl/GlS84riMoM0N9EfEjlMffMgvDdAh1LaiLwUxRjYqp
jrHiR4pUAMpWAx4NMD5tXqMgeYn+TUOtO9uWh4wFpdDGdqhNVwqGqRzrZExXzXw5oF+TfPlikhwc
F3g9+Cykf2ybQKbd15SQDKOPXvTDP9v4eTUqPBwOzT6QA/MUby1VxkofltJlG0s/MyoqadtBuWVh
yYWo7sAUgKRSvzuCI30MgQakkcjLTQKePbViiZZw9bY+87hGL5C9sfjOAF8oNBk0UvxwVnDGf8CG
59TKzMeBAWc/LOBt0gWqYPfEJ8LXOF4DEoL6XeZNKNs4OP+W6Z0bjtP5B4pzLD/E13qghqDLe4rM
VSPV5qYgPgY98+BaRP2GuZy8yBi9xqefxQ7NNtR2NLUDYC4K4XLK8PxIJReF/iHqGzOeXs0Wj5mj
7HDrHJ0PLGE2Vsfl5Zts0oLx7SSP1tDGwfgk+o6jCYMQ3RMlQtR9ZulIbrYDg6J2ixF5ACjCILVa
obcNX3Iif088vIcvANBpKA8rTgdWD3Fc3apOsvU3wEA45oOZ62nr3OrhAxj5fCDLHUnLTgn1Ue8c
vgYMEvI+7Yo0jXbqjloxzwV50rz5TYTOXZ2455npWm0XLFhixeSx3xljIn8o2CSo1fVmbbKc634W
SzqbPAioeysdJq11UDvlWW6zBDSC5wNsqzNi2hqF64L5lsWVwXOG/hABuBYK2DJsl+Ky0hns9sLx
zFd6tO43//9MKJIQf3JLmqinGUnirUpqUMgLbVJ1Ss8Wyw1eWJaX9eg7BsCzN2VrtS2rsQI2T2ky
M+yfzQmhYw8Ln6G5yNPuAkohVe1BxzgGKf+l9r8J+wVv4x5hMKnoiI38TeCUAwUQxfFoP5BRbADc
8od4QBH+l57aG+9faxlEIEW4bJ8F7JRhOczdAdK8exxiiaU0sWZp98sO4HQvcLbIgG5GAMysy6/r
kzXabjVUODcfj/o1DCi7hzzCZNfTgh+mlqFwLE2OaApP6i1nbABPiTBv7nF16mEbLuJ8kwXAckAG
l0O/qYnDE33rqCg+Yra0G0LwcPCcK3yL26DLyDUDTc2qZAikGirtj7PDfhTSXZm1u+sRFHENbJbT
XEY4SYH5npHXoix1S1/liXP4ANAi3NIUSqYtrLNoa9zCYSl5wO0w0mcbBQmRKcLz1lD2WY3g3t1y
DUNeoCpJHmNbOoL9GPpFe5H/oVig4VqfMbAs3tugj4P/WrTB/hug3CTg6Jn4O2itRQAFC+XPbGFK
MmbegEuat/7UnLImMCfYvHr4wbt7wM3E96hHctnIIxJw2FnkiANSzjyJeAV69VAcV5Mei/v9sOq4
cfEI2VTLEMUZK4XWOul8ByHOfybmLzzOybmpz0lBK369sTsvoMX7+1RAa5jgqmoMccKuM360iZAQ
RiEGiV0wc2+mYXST6KamdoKHfDjHSJ0I8THMp2X62YZkjeEL+tRdmMpdmu56O1I1Y2rEDG9+6P2j
jPB4TwPNwS+OqokesCAnuVFP0i2ijYhmYnRP6vN/7G3N/1Fj2uzOlVKiawsBDp8hhjAoQDyNwPU7
NZWY6J3MuGxQJPnRcPs//CMKrp3RfIvgeENWshTbQI2sAlA2xMB4lC7e51XstdLJ52KI8GH9dkUv
pt+DsVbJYmyAuEz867hAIgU2CGUoPrt9QyHgVhrYo6b5lM9FGVRjt0D4NrB77xCSxXFd5GkR1YSF
r68iMApVfbFn+D7rbtAiwtRTuOgybbdBLavobBCQjOvuY4VPRcWnq785c26IBJv083PvIEdX+kLZ
H24xSfNWhOp3Cs43v2vcRphl6W7LMZjl/wKLTdbHwU+E7QTXeFWwvjKx4RUd6v220Khkz8ygWcFL
z5hQ09aveFiZEwc30EGeDy9AZrNvz6/auVBVbBYS2mN29NeZVTpwNuv3oPhhZP9hKrzzynl3B1/z
vd7WPwFauF9QZRsBd59YGNxtctxsKzYMTAc8ak2R3slqIJk8lW2oorgPizPreZ1w4KMmcuZydBIp
72/XwL4GMWzN8pX1NeIHiDmEVt99x4HUhhL6BAUsCeL0S0YMswWh27GNaQC7P863A4IqeVHqgEaU
mWtHcnoBbQWVys9d674Ayef83+u5egGqZ1hA6MyKJoxPpTx4H6Qtv/LrHQeDhwh1IejXpu38Klib
ixlAucMYmMSoPDCpvI6SpIfzyferf0eV0Vm7Yt0U9Uwt0LapRUUERnm4aIKLXZo69IruEdm4OIBI
NwQazUYTDHrXBa+dZGzfBV87MGIjzU0xSf5Ea9kby5vy69hURHJdaGekzeqRgQKR19U33KABNNIc
BXSLHURRdlCntfFf/USuM5YoYyV2tmmMW4O1q+MZUlhuEiyH8TN9EWswbDy6oymqZjfNMjcJzhSx
e4/xmSWZgHSnb/mQ+mvboYMZWCroSKY53l5rowMnpO0cRIomzR5jtXoA8c02ZSwmOIKr+9PiwXUc
oP2NKMWi9OD664gY1bcvvrCHwlJtcKVzXzRB1yYHN+DyXTjuedU+rEcXEMhIYHlv/Mtr+txFSoGp
D1BBIEJy+WelmQ1Fd21XCugYp1/ydrVd9NXIRWvpqmHtsKUJ9tQMiXGCgNFuR2YzYrB7YFRmXP14
rQov4PFNNSwu89ftU8Z/lNb1SDUzu/3pha+IkZMS4ZVRA2Phv8G5Ab7g71yq2P4SZgiOX8Gl/7wn
29Ef2mWBa7fPmMn78HLoiBikYF8fVzjoBjs2Yuqccwd4YnyXmoa9dhNG1h7VylXUteTnk9XHfU1s
ClRAXhZHQT+Cz/JpIFc0VuSbrZMymySqUjlvvPZDLEY8uxM+JwT6Q6dA5+3c3XBHWySDMWoUBJRx
EgjI0ZrCkqISDNF+n9+h/9G9nbRQ/7vWGw7LBb3z/RIFJAFg+Kr82typHdwHMufnu1SJO6dlMOGb
mgOMwLsNuhya3PeBfYohqCxAe3KgOCjigey+ZUraC4csvLfyAkPlSTd5tkKGDUlFjXUqL5lGc5YN
6JBkkuyeyEFqTVt3pb5QnRsYlzA3gqRMGw6xoBngowv0l8WBXsbdvo8Mbouf88nYF0GC2q/BZogL
/5g9IFeZ55C6zoZIQmp8a5MRhDx9flTx+RDHAsulZIfn6p2tFIOwlO1AZs6bWDmLGpqcYl585Hmz
lW0viCNH5JTpqJYhHuMh3OVO493o6dgSbwIMcgSYgcm7AwvAHtx4TQbGsWxK3VkH8ffig4xpB11o
NHjsapRhWsuK8i0ASj1DOB8RjotXyQeF0EybwtZYE9AcfONfoIKfehe18cBZHCUW2gtBpPtkJ4Ue
MVrgBUS8fMn2974jdLvi1qtsEuFeiv6UZXeM0+DNQcFXkLDTTy2XmwgXbUC2g23CKwzZfV9ESuQv
wF68KQ/VoyxAMb5ot8ZuI9o9cCd4hKuxVxuZRasnZrNe2begTkriUH+FZi0zmtt2n9powDRej+32
PW0vdmZQR11UqwOCzQAwFF9wfd7g+SHYCN5VrY4uX/OgjWE7zpfXgpS3WUBDd216eKjB5ETDX216
79Fc6BVxDaPcYJ73doTgQdKXqqhbqosCZ/9ts5BJ5lcUIxyekKrv4AiloAd8Vz3ybl1AGbU94a3U
dyxAo+w2olGA4PA78kJHB+nqo1hUp21IAXGUb6AeiU4VynhzbbFQz64w1+3EuZ04f838+j2dJMSq
Vz2q0GVrsxHNeysJHYzOYJ0UCwi2BP6FU2dkoIXCpuhxkOtzVqffj3MGQzunOtVd44rj2TKFuq+X
uiTp6Dp09ARiAxGnBVVXdg/DzLg4EOehEucFsVDLr7wKm9YT16GUttk2XQRaJkqp1Bu3hrzfgtvZ
h2NLItPG8+3P+M73ImsfLOIBqRrDcsYa6RzCFK3OF19SlqMrDrbCIuWK54vtztrtsMwPqj58mEuz
x2cOmf28K7YisSsp6/fhsOKB8aPPKht56vQcO9Ds/zr3NNk2TRCMQWU6xGzx2ibloSAYJWXvgUrM
KpEx5758ECgDsMUZJy3iJG+UL9fQIAlC5ZOd/SA1Xkj4KanKkWlD7KE9LcBlbF63RjQ3nxEgExsE
DPsY3/Qlzc5lDCAmaRoUGuVtiOxGpITelMkjJSdkZ1rEId2o//7ZxymQEr1ugROXRQU4hE9W8cw9
4eOYJk022tQwWRV1vV2uHIMVtNFEZwnzSIJR7RzrILE1OuyyhUAbqqglYmdLRGWpiXzpMbZRkGiB
9RRUUWw5r7iO1180kZv2lZO3L9y7LCKf0NuyYOqvQInctNpmcXAzr+ZhMTxqJw534LI0umEQqyxI
ITQJpUcYFfbjGKa9wSOM3mBZD4kmjgEkdx5AtRzjMIrtwPWoNQouX1j6XHqqQnhl7ygDetrQ/gGd
S4pG4I+BsyacvcM7mlSrmiEGfzJ0O3MLy8tk7LuNIKC2APAD8NJi6ejHHIkx8kwKwIEZDoS5SDRj
xtJVYFMKdCdnAWYTit5jWIIbKEBsgNgM3FJ+WFuLjFfHQlyiQTYDidi+OIQM8t/Z2XCBd1XCurRd
PRB+ksD8jES0SHQG5nY3bhd4Df9tFrepUeDzS/S/KgiutRzk8Q9Ch9TmI6SxvA+IjJcUn+K6EkM3
Tbqsyew22jARfXgqEeM8y4Jztu6sQBHtFzA8IZ/cxhGGb+VI1QnYSnmIqz8holgbANGV30mcKdem
T+hE1ePWxH2oVCnYsjsLGtkgThBkjPxOrA140SaagfsXWkY2AHwVnF4+MKcoDQ6PzXGt0fwtZ/UP
gBTz8HbsR1/jIZjp5Pag1AfrPp7ZliHxsjjdcWacFhqqtSuEw0APeVfX68pHlriRS1qPeVKXWfm9
/RM7wdJaV4vu6VpBeKMI12pSXO5LFJj2W/qXO1aMzPcKFoViFnuLD+ubIFMjJ5lU39Xq2FTDkgJ2
8Te3+sB7mLDzabDPHQw6GmVyYY6BdMNKn8Fmf/Ntuku1TiN1L6sQ7RVghbExieAybnn5xW12RiYc
j01bMaO/Nea/HmK8dv7uoqB4wjGgeszxFS03e6mLAUn3wYsdK5yXSuDrlCZpU1aDWzh+jaSbHYak
w+DgbEkOLGl+1Fv9YDES1tUiH62SZLhi2MaoFpUqvKANps16Sry9EiiJP8upI5GAE/8bqVOxOZyp
KtXUsxYyBL1igqdUNPh0CbUm30pfdOiwxwxOylRYmeqOdXrj9jFMf+vxZMxyZ9ghcextHKUjjSiW
tSsKxbTJDxv5lDXPcQKFrT2TkZ6xXvsyW0TtqTzUl805bEVxKJReFsTgDsUDYSwBq6c0ZzyEWQ2D
HdG+Kkj1E0t8eB5gPz3o6r/MIVKB4ki8pspZ9nTcc8WWltGLHHArFMsqitk9TXBCJSpCW6FriXoP
rPk40GkSoCWugw+Khsn8pJNHgwSo7J4gvDdDXJi8xsH/ASMq0bUowoxigQYiIVn6d+uzKXYBQBCY
j4f0xU5wo6Sje0CUkegwjGAMaL9oTmfF6gWu8CI5Am34WJ/cKNVe2pmsSGdtN5uXCivk+U2o7rFe
lzwrnTNzYnfNwfAnolqnXCYz7z1o3BMlNg3zFRemMP9Oe92LANVPGsylkyNORQBn0CAvvcMyhURN
FncUYvY9vVYaNbRey2bsij+WVZDMcaKs3FgIV3zbNAZGegYEe4q+Hfibk/MoiMmTSPtD9GbqKeqe
j1pfUrFyiBOhKWAvvoiaCEROQx/z01RW1xnlmDh5ieA4B4oyiK0mt2Xd86HCV4obQVZlYGT2QLLJ
Y9yRUZtiEli5Vtn6o95p+g49RuLbT9nXg6ehS4rmMy9xLlvrUF2lfthNBFnBNHaLW8XJv0Ls5OQt
OahKG9jOlarQ5WHIkjkv4yNYX66hS7vIwCWpf7vnyWtP+am5eHk1z2+9bwVZsnwwO/Qq0rcOkzgI
/jr7WwFX0W4V8kMCqr3kvQCJL94x98yMWdWqHYonxThw70ztQ3aDDow/FCIuZUCnhtheN+pLH45V
0zaHDU/35Ly7srXZswFBRTV5hxQP2QVfLjd1KXCeQalCdYdRgFpMQ5nzMFaCE0jhtEWScFSSTuAY
FkcyxkowPaNz65QVIHVvcBFXfsOG4sLf6bphD09gvXYxhsnZ5fahO+Bxsw3EFxA1ymyOqj8qbQYH
tMynsEK+Zw0HzvAydYwtm/jh2Tsx/D7S/dfF/Rauhn14PL4HkeMI9rvAh6F8gfaHAN1G6XBUb4MH
zG+wqYuLbqTjovrZpjEJR+052aIjBFB943l+hXyZQCbAZ5MDFQfJPQy7abhzNylSAg+EPHc+kc2+
afMZDFo7hqwRKy4nHavGDjw6S/g0QSZyrH6MG4bZ84SV7lp7brcGGdzsyWS9sB6ocxoCRPvY4AQx
2ZnKztBDM6SvVe2xO9t9J4sr7XK6fUFj9n34QZMR8ZvER4kdjDYYZYxcmG9IKxeK10Rn1fQN2HLx
O/sw56f8JZMQe3g5di8VhNjJu8FlI7/DG7PYNCHd6r2TsEMHc3NoLnfnoj9IglOVq5JU3MP1Y8Tb
5vHh7Uj3RQ8NqP5VzdYNCbMV/f2Y25w7xme9VicYvndcMlwimvyf8fLVOyn7t+zqYqffpbkR3JBS
VDAgU5zj9pmuZhQhnxMaAXhjdfra/3dB1LUNbyP+WRpSpWEV2AcyGl2/zYR57ow+CblcLU3GKEIX
rOJpcUE47DiHUG666vqPCwnmDFUe2tdpyb9VOb2Vng08HyGwieMwrWmiNc2KBnO0px+5rhXuzA3a
7/CnbGdvG8Hbg2ea/jub2lPLpf7ODFuz3PLStMQySsah2O6lUhk8cdvacaNpeq+/R3ePG4TwXC13
iwwRWMvoak9Ro3zynsaFkCMVaJ6D4FvJmYXn1y6XJ139Wagz5tWfKzSFv+RjY1oabusC9mxmca7A
zLptFRAtb02zGZDFKqduu40I9N8KNcl1uuCgZHEM/nYTDUyygpicOBlBBfKC1wn8sN7oOHKTQAE5
uOu7RgkMrHZAdetKY6zIIbdByeWmck5CmPOMmXRvWLP5cE/7UO2x3SE8xQCxc65qtxVxqV5CYtIJ
0GBGlwRQE03ShyY2mfrIwuv9uZjtfSOhCR0Cwb9Dq6BRekBpAk5Gb2aqdBTNZhnlNtuT9U0pthrV
ymR0elX0lN9Y8ZPnr4uwUqD5ZoYHFKj+WEoqugcANJnZEjN2KWUQbS9KC/XyfrNDmbVxMNVy50jQ
75+4PHEAJI56/TEI+cKE5PQpAh20Dd/t3P5v+cWpFvQVeYIa2Tgsdcy3zq9DbEIEIXntiaTnGGF2
nOgguc8oYeJQqRDKnyB2CmOPcjU5U7NtY2pvZ/X6d4Z4JozjxdOBdVbXTYd3LtmkmtX7DSYOBbYY
Yn0EOZLRjj63bObhhzulZUf7loriKcMYBisaMa4ll/tp8Q2Fwi6osvCo31ym2xwvu7Kad7ow1hPL
+/CN//axCq2YTXGyIGHUtFcx2US9H23ca+ZZVN2Kx/fs5QaNxiG+0UZSFJ6Onq9nJGQWylKg2LRy
jmwYJS3TlHwpmAgc/K5rHgEsgmVWOrcr1RWyls4ZkBHhnB11vJRQHJBKl5OPhtF9pLB6h6ut4rDS
yaMUNf0PHB8/EBm17dXTRwUHBJOEeWMb1UFTxlE3OBb7HV+V/U9/+r01KNXt4lpEFzHfTaNPu4QV
kclOyuT8aLpoTSocAb+eZPTPu47v7PkP30kSZuvB3Ja1THM1VNdOqGmmm63KZkxGtI9VhePTPWO1
7vOICI3cL/mF8PUEOm55yIA3Vlo+qj2WnOvWh3sruPebRaKK0oA19OalXP5XKeMAl6JaL8oTB0A6
FNLDg41PCpS6vBr5mnaVIen57RzmcBBVO7681SFYK/M5LiLYk0NWWzYSNXDVuD1iACT7BOM8Pv1G
2sPf5uBE+gC6Rh4AKXmc0qKTq2qT68ejF/HIzGc87VDwC9YKxvyEXUoqKKyfoYTUlTMSBI68R8I+
3suYaN2xzLRXBpDLgI9Uu0o0H2LUC/SAe1a6+Fta4Eh1JsfJrRqwTDpNP73PSz40pwdN3W3Qb+zl
XRdiCXk37AUMvxsjA6tEMTqAKyMaeZgiU4iBpwZfBydWaAzzXO2gidDWk4htmoHeXRCRN1TKEIh/
oL1XzQl/MZN3GXnf6J4a+XYZoIZBcIVYa8BCzp9UeQctun3cn9XQiANTxnfNn735zabZVEIKLZcm
mHxub0U/Yx0/pTODaZt83nXeWeJji0uvIvBXxhWFG6OpbdQ8WsjfOnCmPvStXmk4EhLFlJzFS61Z
JC1knT0RQSr6g5z3yLW0LTz6jk6TjUbfVdQG8VrRmqlyLRD+aXk8OXm2i1KPbphLR/ne9OGsjhkK
fobfr0WHTTHCmrUX1D1WrQiRmIOXDo9uRJ4NLRc+zDnTtS8rzZNdMEgVjMBjgupt3LyTi0+twuoF
g+x89CjMb0lEzM95nSd/NW9JYJg86GjWxoRa2OBba9k5doI7v7Mq5xqPfxsrXUAIq2G/GUbcXW3V
WwwpzsrUwFpc/tphTh601bYl+7O32gqDlMRgHOJ7Ci1UIx9gbjAaV19F3Xj2KufmlAN7OnNEBAXn
xrFuCSD6T+80C6tTPq4ZpH0sNg9v8ncSt/lP+1bStvWlgYvbCojPTpdrGOdbNryJ7GLunUdE1GPN
HUXn5BnElZco7H7XR7Oh37W2xgoEq1WaJqQgI4LICerrFOXHES9KldMkWwWi++PYItERKV0wPN6b
51Ke1OAinN3J7OL9unsXf6CVDKxg1oA2U5lCE6lSCY9WKdM/MTCcUw09KtzMRJsnB1YAeJdIhQBf
SvB3nYdmaUpvGSDHqHeeYs1juuLKt+e40bbalGtThTy85KWxezOEKJRhvwVmq4PDHlx9Kkuya24c
lfJ29tfazR8GIwA9TEIuPIuLbtx0z7FfxMavZcEaxZZCSAHphXl0NZWOmLQCPQV0BZ4H0SI6PiJc
+V8watGbl/Xvbo9rvXIjeTdcaTjd4GBI9g/tyoubCQMFsyZHtiFANLObWkU45UBxjgS1IMSqWEHw
AXMpchBtR33f0Q7p2PrqCe9owSt6YRw9d/+eufrcBl1yrgs/6C2KKmw/Iv9JdJE1NBz4sNlYPncR
F0diUD71ZtaifvPlU08pfjUHi7MKPAy8yziKWrMkKYERfStYAWruW+QFoMpisjSF/uBiq7mGF3Zl
ue8qfmlB79svDRo4vGhf64Dsc4LF3heGQSXRmwVrhNCvm4E1TSokQ3vh6eUf2SnEb//datdQfqPC
SeQEzqUkH1b5SD4L1U23WTLEepVTfCoh6/l3d8geZHqugKXbKLuNRiGn19AMUer1TZk7vHkzopOZ
/piQAWDevhVIkGhvv6He36iv0T1BIbCz7P1dBJ40kRnWOOjeekVXitY5puLSv6+kOM6Uneb7d8HP
k0fKct6qgEGmpSqGkdZLN5v/Xib9Veudwpxjzyrqy2vQsHUxVmXmwvUVdLBFLMZ7Vhlef/D3B7b4
QjTHXzLo5rcDhxSen5kV+EfGZpvyrX7snj1pZ3ejV+7LMmLCX1VZbLRqNT1TxxHqaBQfeKbkEvu/
dS5Y10hJRPCKjg/TaEFggehjy30urWWfmM7bPuAyT2WqePrhQmd8nbSpnkf+wRtEN4Myz8HldgLF
ONky2vr+VqQlSC/SuPfcfFRV/i3I260JdIcV7fv29+GovLd0aPQSXWeUlsUQkiUL44fe4FqZCFYa
7amdam0kYgbtti3GcWRwWikTW1MwpS4GCBDuo578BaWWTmxxuESh5h6K2sohOuZ1/7GYCuBFX6d/
+OWOAsSXwHhWCTusCce5OKmOZMA2OV8VcnquLWTrqCG3+fZ4lQTv3mj0ccXD+G6vFxshaEWBrMa/
QaFkA+JT4ZsvKzzsMok6unAtAtCncVADPqS7RCg9yepUWjWdhbTkjgB4bqLZjKtrxFpcy6JQ2Q3z
FYKT/vg5fuGZb2yYOoGT8CADW5U/y7e11qHy8OYj9ovshmdNmaVubh9lb3KqRS+TJB5no4JPhZAd
UQWOB4pqpWRge3XsA46YR3lqiueDe6JUuzsesbxwaMNwvSZbqELocjpZJzmn5c72teR1MewhO4AC
niwJ/KI1wme7nKnlgD4Q6XT//eWFpd+S4up5GItSxojtA11JsC9qybwS+QCmpcddl1qjNsRFGHsq
A3YamvOahORAXu5paUVslnieHhFYMb/hVCov6MC6T7RZ8vMk0/tJwkPnsVuto8HtcJYfAasHUAG4
8leZXekQuVyijwFEXOzMV3WhsaKxk7g/XjGuDY7Pfu7b+7FJpPfZt96xefbEQ4+lpUufejb/QnRB
y3oBaEM76rfHbHoMJKizm6pF285SKBJBM8ewOM9u/zpy8U4+zHK8KrtP8zaqigjyNFDwn2ZcVdi8
/xIvt34BVukqFA+UZPN1y/sfSVWaSunzaXbOX6X+VAprjoo/WjqB/Pi1+b8KIW1vUgXgiVXZSy9o
BKugwUdO4xQoYQ2/MXt0ovo8YiQCkXKEKxn+UfLMJr1lcOvA+JSSaKQntj4EgfE2+IoeMflf2tiS
2Bb7PLo6fesLoB7x1WXYF+BW9IhsJ33jsWjdPnsLkhZeKHgyANu8pwFXWjjnmSVxgtmakxlmaAXq
1R2Xbe3LS5gXW2z8c9UpHNWQ7rjCUlHp/0+mm5PjbGuhyVbX7KbezjRK7TGqKKFNCMekEiAdwRez
nh5CPzvmZFKMP5x5uuCS7EwW1TH5dKbwAlacOXTpryyfdp7QI7KYpVakMAOVHwhETIDr142zAT4j
18fUIzq2oU4COxruofBv/g8xi799RuY57tJhTwt1QobeFb1OteG3vCJiuRjDHrQBw7cG7xRU3VuP
9fQ4X8f7L+wMfmHtVEk1oUOyERhouRMPz096zTPvou1kE4bD0cmoyV+e5O/KnWyEJCSw5pqUYg39
wyCI3+1SfBHQ8s9l2hdX7YoYdF9i4SW4D4yM7nv0us62OtKpP72erHRfqiR/RYBPcwMfVEFwmVJO
psMWyItHOuBYDP7M2gXtRem87SgNQ9Js0DhYjpS+qW9iST0/3ZPp4Yhywe3uobhUEuetToaYDKHD
qSULul2gdIsI8fy6iyBFrYjeJ3wtNZ/50ev0ZDUmfS88Cl0JRe9FBvXIRbf0rwuYospQTMnwLgYS
i2c40fLbJJv619YHWxv69IqQiIgxU2ck7otxjlUWtn9IXYKpennjZyWQYAs6yz0qfR0zSH3gEXXc
SfHGQK22LJasJIkWxZE3LdZnOcPE+DTXoRbgzGcAzjcY3QqL8foTPjUwS2UQJAM9BVmbq9gFKM4/
4GYFP97QzgnkfQ1Z8xlztG6I1yxDHPi2XBMWcRNGCcGOOeijM3y7gftq9jZFO030zfkKGMuN3Fd8
Uic0+1J5gX8i//B5L+RFZKjTC/EAhglagjrOvsq5JW5w/QdwryxE3sXMVX/p642bWffO9ETsSKIv
F4jfQ7vbtBOwIyTK+/E2/Om9WIfyCndMQC4Y9T3XdgYvUQvJOfWblE/lPzSxsO8J8sYupAO+y2kA
Q9igmm+k+aF1BiAreADuPhFk8vaDKC1FzhtBZM41LUkIqNPvjkfeObQJJLK5P2/8/xxIrZ70dy7O
UBPwp3q4OqqFS+DnLQov1ux+QFzrfb/ZlmSYBfVctmYP+My3LoXHQQ5xRpKxB1b/Bn5nGIWhCWkS
Gn6OgKzykBwNWxtbr702SBC/GU1QoEAYONb+7L7E3JdJokUSNObDtU0hCYh0AGyTGYK0OzX6sQkN
WO0qvCb+YK+2BUsIHHhRNZOOpTh9BkMlVgUJmF9XWux98g88hh9X9zp1fRfCfOuO4yG3IFD9efHo
xTVYPwcJuz3izjp7VS9FE8i/3wzLSnzvMbI2fQnJk1+zYOV0QDy5cR2hTHisBzTpTB42c36Fttrw
h1V+0ceoQACM4zITyO1T8rMI9YoFMqt/N4BeGHMUp9BbsddhPT0QG8wybJzTJRt9uP6/3b2K8DP2
RQ2HIpywhN7nkduJAWim8Lfh4JMzYLZ0pXE6bLA9EJeWYSe4tkNJzOm0CpUZOpCGMkRCDc/4916w
pzLInIUaRSlB7UmE6pE4/vihKp6psQaSy+EJB3Lsm6HmBKylPT/N6cyg+bOgX/DwaTxp4KveCg1B
H2AJGsNR76EnoYBRr9OwaaWrhkz3JEHVPRoNRDFaV2sglJ2SnDZYntfCtnrmosOO2wtnccRy0LYk
7iXhUEv4qjQQaTvSPgDtDtOxcY+oV+KsHjOa7girNOIwNMLA1inNkwRNp8PXzCyN/1AtemhpzfHU
lyH/O0WHjL5s+bo3d61ag0CnwQ6l/xx8ygTJ3ziX8zyjUDVlhx2YNuJoyzLvQ89CTI1J+7vwIcD4
9Cl0UprwBItaRMMfS7qOHnt434qWJm+svlfJUCzMUPX7/x2j8qCTH8lg//HMdo03SZ/5RXGKTw5G
K7VzidUfnSw2N6+UMdsX8FLsndiXDQRPdyJWmlwwrXRT+cBf2LYx7SGlzN9RIGxC6bX3SeHLkyaP
vdQjaZWLx92gqp0cqu73132XegNTzngcAJo2aCR1I5ExAZUWM4doCWVhMzM4ZpCifUTwQ+7+Gy9p
0uB8g0aBR2+RZ8DFGWwuOEFHtq2u2DPXAeAColv8Bp7OUYFDr4YEWJhfO4CIuYhs+J3ueDYEGfz5
E6hAA4VwJj87/6FKtO6QeFSLd/2DxXJwBSjy0bsl+E5kf0KHhkzsddlilpeYbY8q435kaYiQvYok
hcIou8l5c0784OG5KcZvIvRX7UeQDnqunV104yQlpCI9vzAQ8uQdmG1S+VmC+pr366wo21kAbr1p
yIlBb/aCdM5hFDoWo5md4G7dzJhuGbMpOw7j9Fux8Dnmc8TQD0a+Y+5CnHJ3KrUILellh9Y+Kt2M
0LH2QdHvdXV8HoGhKPZx+ZmudHn6ks0H/NopnYt27QeKZfqbTNHLqR3MeatKj2GHv9At6G601Z+v
RrI/eAbuW+SYUXZ4x/DKLDKOam1hwgh7ngWAkvOqA+4OMbjP8QgLE47FS3Z59yXVtABFmTFvQPx6
1J+wA2iQsrg8zioZC96cxUxUnONA30Mh8gRRWsMhICPI2QznAx4A3OiQ6axcBRY488/Nlrw9n3Ug
06j+k9YnXk6ORzDolwRR7d0V6FQnLnOVU1ZZw65rOEMp9l9O2K69T/ZIDeFRX4RcxjazxJl3hlmK
1Jgyc7QkAOZQk+l70Jv585UY5MjyLhyrkWLlzM7bjKvSfZxcQ3yeLjqrH4XyK10LnL8Dssf83l/1
lU+Qazq3zvR/jZr0xSzP/nw+1rcGg4P+jKCLuFTLay31zm4OYbQBhdeo02CYX5D7Rl0iiAjciqoE
z8CgFfaIksPSxThzqFnj+AO6UIWEQ4PlnsJ+pTV+1jtRL62jOgEV5eLFtpbQzc9FfNTKPaR83XLz
wxi/ClJfYtcdfbuqZJx74HlCylRc8Ktak5xvDHP+eXYy01rZFH69KsqmCnSpWzORGoLynieyeSgK
liMxwtaso6lJ3ja0jr6L1Pjnwl8d6bnaqOy0qYzegORKOFxhAiL1Pejr9Fzo9dsNKGW9HWPdmHSD
rvSHMgicQYp6ZDWqCTaQ38fTekTguNHme7FWmOGtEjFlLnxmWFh7CWS2vNgeMDU5jWPYoRc+JCdl
yiJqgmNkOL1gIW6FxcLJmNhxtCJDnauOhg7P5fzBTyXrDPmEv1yvxeWQoBhGbb8nY5Ane3UHp7/J
bUd2NNKW353P1+wnGMKuA81NvuVI31b0ipZqj9Pe6qEBpSz/NAP771GU7ynRaBhd4H/MCyqK8r9o
l1L467hNZApE6tv8AOtXrNy4yYaMcIF2Kw2UYdK30h593y7ox8MJAxm6ZNfA8LFI6DXotnWY0nQN
0NeuYrYfZAuh/dSmK4UEMyJztgHuIPVWZhcDwxyKxFDYfgC0z9aQeV5znhVg+8HvztObqqjypnk0
26puN+Kl4fFiDR3DEYzSzHnehkQC2pfEgke6VGEzMRNHyY7kpnHkwJ9W0zm1O4hYGN0siO0KrO4q
LgeFHhrmrmUkSjLBHbwQRn0s7sVsmEKHqaESlC8fyxL8Z6Twa+u+XM/6vGtrOc8upLG9kvuXGnfU
A/H0g7O4AkD1pQDtk2X7OCIoLvFPSy0eGxFrUBYxVJV6aiIHxM9B7OYE3LZYBmYISlOcnstzenrI
WZ8H9RPYBA9xjbq2F58gSIyufHgDR1E0uUzaa6KWC3S1ByLvzt3q2n7WoIdtsHkeoFgi4PwwvPv6
061ciDJnhVsZfceHvNTkQfFNuOphSLhIckbJBcNOIql4JISGtfzIYHUiGpyH27fAkNnraE+bxceu
9spEPA3OP6YhhbXdr8wI0WNNQMF2oiPfLy4gHSV9Nm1MlX7QcjOXG5+WFCCU+KwXh8dHu0lEQ0bA
zy72+3vFcOAxiiQdfMcisu/ZYxlo9G4dZ3QDudGM9oAVYOWhVRHxMmVHjT0dPcjrG7hb7Jx/l/NF
EN4Xa51Zq4KVTbDysIghHO/3VE32CQgbt6AkFrCceT1RVxp0GBdyIa/MTwQ3n0+X9ioReJcgkkUh
F5AKAWZUd5jwIKOP2PZ2C90KGP23OmWHO1F7rsMJ/zkxxw4rGk6o2V3W31+0eTGIts8EKqmel3mg
QgphBpRhBF2KRU/Ez2U+gCuFgUPTm6/XoCAGJDyXYMUB8oC/8N3B42amVtK2xCSBkLNMPGba2Rib
jXqYdsQotu/i4NdVlI9URCu7Ad38+nCpaYQvF+vH5j8et5IG1t6VeHItWyvK8KCxol5E4zmZ7MFK
LCdA8t8IsnIHZ6WhxhgxjYjxA+ks6lmj/pWJkI+C0IYEAkvOuRClVUYonT/IywNFP8JTigFFxujb
PTiSAoACCkDEfgNy1ll2o4EE4glE/CNMnIz66jsUePToIiJ058bwN1QIPSk+O+yrJQbtb/RC2ZbI
5z/Q6Iyf8H/Xt5g8XBSy44xj4t7yA0QKWySPyCpSNd0NEtYNEqCcfYAYQkngmfF+8iUpmKTSAfjK
r4PNf9k5Jp/Cevhca/mSf6pFJtG9/jazXKTsJsA57drhmsipIYXEHtQBS1Wyni5dg0/+PNjGcNkd
AyzT72xSbAd8XtmzJvslnWjQ5LOo0I/ymjkcCqOUqZrLE3J3Ibb/PMUzZGm0yEsB2m/0zJ6kFF+L
UAZ5mzdAGzl+0pMayqoLQJ+G7NeDzk4E/5Ecd8MQaMrYZGCK+LPAzPQxrxQ/S7l87Q0sN+tSX2JN
cyc/n9kxyVLrOD5uLo7JS1CedMAqLR9GNB2GNY6yKy3eXH21r1r1BUZb8vxtrpzGJwAyHbR8J1k1
IXgHKwf0xjY6XM+wdmwHlCXQ9KvXM2y4757Dqz67HpToonRbCOe5BGj0j9QSJbkyv0nZu/stsWhM
fmtFLgHsyVMWwYvd16tk3ZGsC1ihN2HAY/ml2Mpubs6H4JdNkKtvp7zLaky/YbQGnbun3Pr9tzHV
fvze0oJ376lh3YZ4b1PBfkSCNZGH2E6EeTXJh1kJoLoZOgbhOvtH7n92rxGCmlMzdfti3/zv5+IT
bZADOuuZYuNnOxotXIgx0O+ORpYKIU/e/s9Yq7U4bXwCb7sl74tRjEWd+QPLxyuVmMYipz3XvEPq
24hLSVXl2QnAocOfg1TQ1wNFsTwdZWGIDiZ0IL/O3QAMBMlWeXLYJYOnLQV6fCXf9PCHmg95zGZW
GvLeY95pFOwmU+6F6tCOhGORlwaAVuENXL/VpfrEnME9RuK4pGTJ+OHOKrAoxnFtJdRDxBhppcTc
IVuz25Qm4LwXejc0qCyQNSNSeqv/D2Q8qbyi1oeGXyD9skOAuZOTW6PR8f2l+ISxTpBtS2eV57us
JuXHw1jia6UauKUD1atfFuAhLs7G2PCwp5cWECXWU71cyQGoov6oDCsyYlmQ3F3Tl2K0sIT7RPsu
+7eKgU5yZbB3NUlBUYdYKY0EZ08ZSfY3RuwMDL+oy6b9lIhRCPvlAnHrfFyO0VbcZ5Rdd84lUFLt
9lVZBRtIiTjYkCuqxZ8kpa2jOPG3vAVovO9JvFR+vlg15sH4uDVmAGDXND6PyvUurXswoVKekTl1
QrZ+6zxaPDHiEBsUBC0CMnuQmC3aW8PSE6+pWkw+9q+YNr2dOnA/f87+M/DJbFtyCdvAIx6fTzOr
Mk6b8e3Y0Xi/dPR5vdGlD5lBcBfTPkB1nOsYLsbT5XkC+4gGxDxgLjWcvJIiXS0QlOk3ORw0j48X
CLNXRr1Mx1X598wDAFGB8pXpNjP68fa35jKsiUG6ZrLsymNo0IJ29UMX5D4dPwwpAY0XgIGT0Rfz
Y32EEVlFRud7nHHeAmZm985AEabKdrO5sazMm0qcOrGVYB5Wg5GUv9T6ZRAPtovoNZdCdyTVeplY
vVJz2/YjEuBjDsa0DWbHvDR+O+dQ/QiEa4V9hAmX28OiVL4G3/EEnMLjtaHrwrvFFKt3cKN4KCw9
YnJ8mf5RGSWOe8cvS7A59yzrQkOdOFiKt8phd3Ztt04H5LUFI8khffGbwwa5ud3K1p8DRrDDu7lZ
DSDLd5Cpp1oVoqQ71BGD0oSswhooGJU5+lhXkhy7FEWJhtS7RbAve3z5DezIoFhL40E9Edu1Cigg
mzR/e28+O9PQiMIOjH33eDYgqcCKkvqdhUvI6n0Us2omxeUjcwqHaf3wAe874Fap5XaZQxelI9V6
y0Ri1ZjQGkW+xcDm+kxkY4GCmkV0s0yi175ZGaqIxl06dhXAgd29DrlxBuUngAUaSMjewweOgjLU
EK6XebYV+SnFkf+4J0L7/Tl00OmifzefOtqBU5oBWIRXx5RUYQXis+edhCMSYyBfZ1vl5AWtTvY8
JEMqfMeGk9McjriK2XH/aZwGp/WCZncD/+tULzcx/N3vzBAXDUXy52GMyygLqEKiXG4j67VzJWJg
B2Opsa81JSVf/ehJ/NUxuTh1iwKqvYhpavdCHZ0A7yccQIBxTbwTX6Wg56oHfvov5vVKdCrpyTmn
TyW18VJiIPgm6pheEKIHht+Q8q+yqNZTOWTFNWabvXDqjOjDVJtBcOupQrqVwD/Xnj+ZjxYFBNiY
XKc6kV3g3FIA11q4BMrBPHBpnicGyJAlI8pSbOVYEEoWWVIRCZpwrV7ahcQR0YQcYtF+e1Xv3VIv
WKo5fv3bw2hQaWi/oOD74PAXcAyAMnpR8AjU1LmjRDEZCBWUgm9QthHNoAiuH6x+65JSKLFZKZ+s
pfLLJ4rKYkuanUSzqIHkmJ7NeYBM1UFD6lua2e00VM8lUPqKWPPZURjIPSDEbJFXk2c04++WlyYP
9rgGNNk5b01whoaD9mc/NJhbh/FaS4zN/z52nn9seBd3OPH/gwmHwKCHEKyJtdx8krbWFfGdBKAn
/5w0ff5PY/lBB0gcfXtvxOQPYJQVME0Kz3rwWKdb9VgkILqMeiKecK3TyTJp58t3xmYsZMXJtQp/
RCFtxuR/E25A6niPwYOLko0Oi768U621YATZfuz0a+USJY7bnStVVfXBoCZLH6df1f1yx3KI+CBN
K+iXOiBWfb+Dea96dck4TS/7J9y77BgJaOnk6rJ3HoLUU7k2UqnnpTkgWWD97Yc2veN8dURNF6mK
OITovXbRjefCFAvjeZJCHLxRHNGXG4bF8zcA7rA+7zoIMy6/f8lgzdGGr9/EmoElt//60mrDdNPT
lRNDqcnM/8ePGeaKwRSAcSnQCiQ4QCz3ALsCkNAFgAP9vLmyOXNuMLQiaoZB9LOKmzt4238hx95+
NCRwUm1X04fsPC5FVdWw5o25gGinEaM+ssmVTnTrWob8p8XVO8lQDoPAwnuCShE7uEHFhTfQXk8z
pl6YGePZIckyNN/pwBqlQGXCpyshl6llKwCo6XwuMu+BQQ4RhYc4y9mlpbDzxpEkfFcd/kQzfha8
X9+MNqu3XHzce8VYXoUkkNYJ9LX4ZV1N6AyPtx/olnaU3Q0LmORDPWHSZRyCT9AvRysX3ZVPV5Gf
xe8MmDMbL9T/YQfktORImTee1a++JA3fihmojaM0lWhO/Fe16PiIKWySN+PXMQLrqw8RzjGaC95S
9H5lrKjPk/xCl3L02BnaTKrLzGY+9/TfbNj8ji/57MfES3JibcXQg/5aWjHx4MxANBkRB4FEHTUV
KDHTxPIUzeV6bkNiJhRvQx38VftMu66H3pffbIlCHlDCkIOsMggSU6R9aI7BZg4S9QTAxiSduBWV
y1rPq4SbB25UEhGmq0vs6cPG+ycQdKFinm2U/G2RuVCUyIyWOIi5SdH2mzCX90rNrWzVd8VHkYyy
C13CPwixP280hqZDtebX7qP4SknHYRWvepFE0e2e7pvDgY6Zsph2kHxKC2FvtykHJPPk1AIQ+fah
N5WNo+SL6etRxaYvE+xPq00sF1LS3pCzxW48hWCG8hqwjOshm3DdSnCmcWKTcvaf8w1wZhiNHplS
7cBKLO6HGytlH7L5eFDoXmGKHZHtDcSAUpZHNKgoSNu1fPAiE6A/XWV7OHMZfseA2UV+s60PT3La
UVF6Z1cinZwY7fHcnil5D73aABt07p2dpmhmFQ7oGp5GXOf8JraeMoIEsNZ2HEvwDGH21VYTOjvR
jFB2ZaZDEuQdRT+aJjxacYuyi1+992Wcy+qSBx0QVZLf/qS25Fektu9JIg+oa2dASsoqAyveY5AF
ctUnS2WlGCsWtb1L+bTBDgMuHsdnJi3aRVC3VIx4LfvNBZvYZn+dJIUYeY0Cc1a5sIb/NvUS2lEn
2/kWFKclcXxD77VzcrecjXAgT9KSwd8qhF/Ja3bQRtnjJ+iWD2dfIM2QqtkRlW/FtgT+vybvkPel
FBocWaGnYPlbvFs1OYon50ChvMOtAg1fIt2Z4P/AETOsklrT2gzt+dWAko9aF8wpHuc89iJ3KWU0
IP1IN1OsbI7Owq7XSSGvDn5wshlkx6ZWcgVZ5GzaQjAs8yWRbppEkIUdwCWwtHnklRYlKB6/OvPl
1JsURlQDQcqNyOWypfKQg3G9X6IbVZO2RwM0zWV+7UzvG2lkiXXtCyjzYRcVreZgBZFzGNliP5mS
4qSEFyC6kGSYkTvfdM+5QkCHoVWjeaPyDh5RliZY7XOjZzdf6ZSitYYUw9pcGZD8smDD8QaBMuHC
xUGLEC4KefvvmmIMI3RNzgppWZkhAjNcJJU2CSUb2Xx1khPnbeaEeq0+YIpopR4xMtbllJIpd5+x
WwZbSzRtK5X901FvvRKCvhwPeq5PhH5YGdsBwAyragWObwgnBE9mlUEw/49ib1er2o6x48zT1fMD
5hLciZQ41lu7nE0IpMRwg/S9D/QLd76KMoUcjClraqA0KSWwJptIkSbpVKySeN2YNUcrVQnyVipE
4z+bQYumb8ef86FFeThVk+8d20G3Vk145mFaqh1p+klTeKxqUmU13lKeJU7Xl9hbIJMX7Oq/iANH
r+sBUSJ0/oEHfjRInBskC6r8te4rcXXQpcRSB4WN6RXpBEjk3Oan49zYansBteW0yIfwUtMai0nu
mUsIQpYWIfviWQHtVL3+Ds8n10OdeJozm29F/mmBW0789lRGcUlbF6ubfcw3GtCuBdkcBmInWJ1I
DYNZITYrNhqsra62Dnd1/d3p6vc/k78uWd6GIX6IFfW74wnets7IDsSGjkJPfy6lLYJi94cN8cJj
k1amhQfIqgO7jYTPzsCHrgKh9hVxo2xzRuoW4S00brJ0HC/woIZHjxD45/J9VtWs47GvuIJ9zz8S
zjSa1NRMa8X4ECktto1scOTHzIhvHI8l7GG7M99nRicYYSZu3I9CNeYzk/fR+w/+bUDfQfTvgETc
veQX6EOJAC7F/3Pzh3jkBbqDgDOIXZ55XV5GuUTlU8S+TpETbGlBGSIWtc73j9hErG41edkTeuu0
RfZ3pvjsp+PNz0Roso35kUf+4DLBZ5SW7/wE8hV9FcHhjUzwE6wGYNR5Oz8h/SBjJbfning9aJIf
Mxu8oE/oXStVAvCxg/VZLrIhza19rhN9T7r0Qaff9WOewc9HuOumVBlJIQ+b7ECXKCXE5mI+FCOO
pHhI80WqBppOvhftIqU6UDt8sZqUb8cFYpYzIc8x7ZGZP91LU1lOKVK8ZV52YJWsYi1jXhORQ7qL
6dSq1F1neGFD945b8Wf+LDFhKiCF/OntndbOwjm6XejvVZX9lQpkpGx198qp0o1uYXrSyuNMWYmn
fqG/Sxw3npbCzbo95ASPOo/anfl4UWxIk/ho2hKPNtR/jbOZn8fCf2+yOcOHU+fKfMI2TFEol8X5
5RYtW3rjwCaMTB/Nv09nsu23SBrewZttuyioXxyA2R7QdnRCA/FYh3mwyPfMCnfWSdzFED+Y9gXD
jOZw5lrKZ1nd/wRVwiUrsJedZ6XdA+HXcKfMtTI61is3fEgDNxGp1jmw64ul3Sv/inFA7EVzD9JT
rNTatfpjmQN+3lLDNWcue4k5c/sRxRaYDY0d7GtqAADcw906noUHeZF//60U0QKipt7RIF5i37ds
ddQ/hlESgkUCKPIikNMDIGLrvrTdHamuXm14cpI7nlV+pkb1q0+N/it/R6RxShCGsCzfMekIirhM
VUjtVfHpQRMqE2j+YLqXoZ5TjWDkymiW366w6v8U5Szi9jYdfew/hg/KKYdHQxVlZWBTdmzjSzjl
I32WuWTq0PUF6zHuucu8M+n6O3yJULXQr6jlAQCAXYODCOtU2c0QC5LH2YpnEy5xfj6jBnLLNeLb
q3h+3AsFGKwTm246NkFpS78O+hhuZW8zIgKoyraXPb+qXPODjiMJK6gs7skBGGaBomxzK7IqpLVG
TupRMSShSm5nZsrI3HIxqq1eORzCvoOIARXRZ18v91DcNFjrGxldy8uMCvabDxNlWNFN87CpKbs/
Odymy3GiPe9ITWJUMVwbMSZ7G8QYzN4Cib8Vp0gxFuvIltg+ZvYrDX7yigyG1ejJ8tD1YwKi7vg/
BZXjABf3R36HY9Eg9jNpJ9RVn+vGVb2bnHv5oMdQfIv1RhGdOxD4rAThphevV4MyVxPno37TddEz
wZeIsGGi4tZBssGTbgX4cw6oXaqfqFH1h/CLJQR2b3qnXV9limxPFCrzFCaX0YaJBb+6tLp3chxD
qNK1eU0PeYPNHhK/UOPVOHc9F+5TSRiwAC8qbdIFNt0hedwnu8HFShXs5bnbCt7LTSlMfWc+icGw
EYPZl7GXBR1vjyyFm0M6WfYLTszzilUbQubhKw8iA9FJ2nJ//Q8YsBmWRAEJuTrWlQjGs0Iel6mW
NEH45ym3YJAeFeX241vxwEa1rQg8pWX5X35ZgKP98TrGCnSWT02XI8Vfb4FMzA01Bgf6NQNA5fGy
8DwISwLtqjm8OSUeOzTjwVYHa8L3Ezde4iG27jYdkGcTGuIev9m2ix4Xac+pXq9ZXGNX2MQuMmax
YdTUfRSwbtTOQUNgsn/1JPWzpERVmrWVLSvhYSPP2wxb4OGrEIsdEioEHBGkcWUSTdYYArPxxcAc
4hJGzJrARII6Vxf9AME9Bdg8YLHyPQ6z29CqzgyMIimkGiN5CPjCsgEW+GCOYW+JnD/jlWtV1VEt
BD8Ej9lLQBQC0crCn7fk7PpFjt3C9lKqBs5X/cL59sSuH7Gb7DvkYDBRz0BuLYJheaHcdxQUvLTd
duLVDz2SkrfYjqdrpWcUpxgSc2gbuwU06AP/l5IhPs9SbXDKVOMT+bSfrAYDmk8fkxUYqmNYyCtQ
Zl6lMYC4AeQsw8SHjR8TDfVHVLzp4H5gG5vqrQIgLwmWY587cR204kmTbj1mnaWhT4n3NBOMLiqL
VlzL4rg03an0yUCSydY6lGlt+HzqyIxXCoRnJRNSI/SFlkh9NXBaASp3X5zIqn3m9Q8Kdhx0JfOt
2AL55DZursgkKWi9u0ZszxkKaq266EBBrmoPrGtouZ0nVuRUOs6/rAn6XVjpXdGGZe6t+2tDa7d1
kiO8FCgz7o1sXstKJ24fobOcNAQAV/0K4AzmH2LBEAwbzjsNmDJuybpqohG+bn1a62zIgevSOJXn
mR0AUvkBzpwFidLmP02nVvfWLzgOE339+XM/CRsDfT0vLPN7AUdqGZFulJpk6Exr+qOvUSNWEq71
i/DDQXmYh8l7NcqxvrbMsBRh9VvnwLkpKdjUig6ofzaa4tEUt3GDEylm13gRcN0Tp8jLE49y/3b0
RNLtxcbMF4c3E0ssGu7I94UF+Gm1fvAi5n5CFLkLap5BWZ/gNSCBu8cmafqh7DmDVXvSk5Paa6uE
BqIbHnE/79VpBsBEclFGTMNcx1so3Wl+fjH/b+CrAeXiXNJbBTAdXOy8U9OIqeMbyR5Zfbh7bNj3
mGBeviaKUmDNQtpgmMvAdtPkkmRC6I5GhCvIklEUozrGo32iMi34xjs+DpZ1CeiUeDaWBcUq/GSt
vvriP6HHQg8OFdOiABhdtF18slo1PihRTgKKOwtFSjP6TS1wGBea9vkQcP/XRxv+8izCFktjzI14
6f709nGGRqNK5v1lV54Y+ctb5/tr+CpTLuScTAkrLM/NeYGykldp1H0/TyDyYmS9KiwWb0+GhZy8
MSSHP5eIFPnwm/V0cEwnYNcFigAATiRCVx5acyF3jRkHAE7IFlIXvkfZI0G9CsMm40Us73BTMZcT
cNI/N5mohWjVZXnqSQ0RXzRsWT4krnM1PyV2k7pxaO+ixM6l9D49os08OXgfcIM1nJpg5WxqYK0y
ceKL3cRwMCSm7zq4nGgmnKmzfBE1+wWVYa8FIVInGCOeMoXLVJOb64wvVgeQDnoO29X8tz7Q1vpx
fq0SAekgShN0Gg9PI2FtZ4Lz6pXAcfWwf6v3BYttV7+mc0RKOTGA0WYa7kj7G0PcOjk4xpCWxiZK
KgyuKhalEtDukkaOmYe68eCWjn6LPvs+Dkecc8DY3DuZWxwW0WW1Cd7nE+ZNz/QVLahPbFX3B660
E90mfV68LhUkdY4g5gg+xQFzlFV23TljwmOYp+HVMUWyK5XQWf/APFGIX53OJUIS72i+ETbmp/gB
llrfkbS8aGxKu5smrfoOGdIu/UILUb6naip5xMwVUdpjvFSGY1ONT9j6VNmRAaPsnfo7DB78QoBL
tnS4xoDEWvH4m3HY2GMKJEzedp4IsPmRUyyMHynlBWbPtabD8lUtOA4LhxTbe1/NsiMhQT8Kr2fk
60+C+Ef5Vm+CohvJMiGPxKva3igggfRc6odVw3Kbj+WSmpqflrTImDBRegelVUpinL01eXGf6v4l
t/cnyLv1kPV4FixTSbHXJ8rrcizdmS/J08RESYvfddZ2EWFbT8lxm0cMW51isQP9OXJcYGtQbtbm
ecDvYI7RHiX7u3VdImxvOP4fHINJf8xPEpbzwYdSo/p3J8mzSTPn4CcLw7axRLdgY8PiR2qr6eZh
KLTOkxXCWPWl5pP5ZP9ZTqkKT4CddK1h+kIhiQOu++U9/LeH0j/EXJ7ErFMqzqp2z7qoRfgJCzYU
D+35t7jF5zPb+CpLilCN2exLQyNECcZ8rabbfncHldZFkGfZtWnHMEi1MW55JwPtQbnsJdLgoPL3
JD21D/d1iKHWPvTuUZI4yCp4WW+q75/AACKlLlElBL9IAtF4ZuFZbxoC1U3P1u/bRjG5/B4IXwmj
sVlNajrrV1UtQe8JssJABOHirDptCr6Xj6OA6NQ73/uhBvsv6lUa24ZkVibi7SjQq+OBuR08+CG5
tqp7IEhiLp5HjvNZc72emJXgT1yuatviTslZNdyYeIvuPbDGwGzWXliPUcv6rRCB4OBg/Yy8WPO9
b1J/LOa2gvaDAWALqkuipt3ZfvB0E2RNuatJvs1oDh2di/iJXZ42mB33y5xyhn0vv29EAd8+/eoZ
CLpWWoHDDbrMQNP9I3wc1pzsTXHoe54sxEWrIuVHa19xTZlFlpur3rT0Vmt8Y+i34YLqQ+uPFgBa
iV2uSraXr9hTRwSBP0zKnd65Qlg2/NsiZ7B6mroaIVRkOgaavJb4kxp85BVSmGT7BUdS2uhKcY0O
UqGtLZMaO6qtFV6bfFyy13DX43sWMdghVMwVDt9W6Ndj9DkSc4SV3g257ZwOkk7YFzESJ7gLelYv
Lu0pKimwVEqUUQDih4jAofjLUphrqzJ8SvlXFFaOERzIdfglUUMKZeHQp1MMZmF1jRrJrNYA4sWP
N3WdeMlt8awUXShWtsq1wuUevo9qupohqhjigWNSah+2XoPt7NtvhSMk1IWQ3iMeXRpevcz4Vhb9
DsTUxuKwd0aHns5bI7Ob14HOGGSLsMpW/5w2Kxxe5nIUFyV+e8j4DEscWpMU7StT/xW8RDl6q8fF
xndu6LvAcLoQ23g+qEO+mXK4KIZa9DGG0nd7vJl90j4jmP747GEB1PhLraw3XO6WnmL6KnRPoJew
xYDSPmHXI5G90r84sL+vSi9pvIiRmbOfmo8ZxQ2TP64lL1Yn6+Pdekcc+P+KqnvO01iBRRq5bS7w
mGX/hDhP3Ky21qYzZ80vH1A2WHmwVxfdK76YvJZjN4uZGwI2orWAB9eaZVtY8ai8bFfsklMk0WUx
/c3GrOQ3BemO9j/1msdGKGPfZ67MJ8YYoyzHgq+bZo/RNNFzoyZAG5jzYAl5B7TDrEXGFlUCZhtA
LPpArLG5gw42Gv0yb4IAKxwIqI1K9Mw+xy8+vLc7U/w6kMSkLZh8PE8LHT9JXqLntxG6DLPdui8L
gWZbuC90pEdAv560z+64nNIPZkC7dBJmpkABM4iwIlp8oHwUAyANE0tb+7J1ADmFWk5cdJJcJ/CS
E/qc9d6cvy7J4WhKaKU9bbxeY6FXjPI057WMYGNwu6H6uZtZmpedScPh3KcCTKuu2z5sejTpts72
2jg8WHfiD6aMUMGOvZrm4WFVmdF7iHQsLe3/QovSqotQQFH/mmEUD0gNLbDdosgEL3jmjvIOtEta
cd7E76GMYhrS7PCkJ9AZ3JIJlrX+aD1Nbd+b+QQN7dpqwZxidr7yqT/6PN7ElacBRjmJNk5Mm8JD
iqlgNvyE7n5Ci6SirLjfoBJ6jh2EM5gP9fgSaXwcHmNZpmGFXb2R79F9wgqaE2nLCvhuTT85b4oS
Y2Zojmi2ATpwd02zaYfieOUzvb0pLgd9LaxhPxQUdsqqjw9Co1HpON/5o6hOPnAO1nExM4CvCZbe
bDEc7nQr0YT+UPvDHscTkWiO4umGJLMz/+RbtcMCN9MTjK7c4I3LyyB+eht8F9n6nEN25+kFWwBv
SjEKF/AFlm6+PrVz5xmuIImO/W5GYRGYnfAEEXQ5Cwy5u0ZALYsKn3ahNXYqXGRCZJn4Ai4dwt9i
ileCh05bX5mkYTBLsMO9trZyF/YTsOg9Yo0kxv8WUCZaF6qGoT8ew4Vr5MefKtCTYXB5hc6lQNFc
yjaxjKPh1IFFV/Wbg4bDzNOnmA7n0vNLGDS7+oyySQT4JAd2/9BG1UkuF5o4yYb59xXGdXTaHMLz
IYx6M6c3LTsHJqVMmzzszUFQnC+Q/ifbZeBDo52EtbkH7490gnKI8Rs60KDWYekkNyUg+hoGeZxH
XhyzJGXRgHQcKa7v+64rbwiQ/fJPnzgXuPoP3TEiBdliJbA67E8AbVnZm/EWTYON56s8Y4ymItIc
IMaaqjBZrRNiFCn5QGiz+LhwsdDdKHMmw0rPQfBrZtS6S3WLJQqYFurzYe2eXJKkWeV0XWOVwK/d
hSOZp4FdyO2o7gwQYg+wpvFZsmoNlq58aVt2L0hBk/qNbnTyFmVhMZZZCE1ukkOvRiwtrXkbRCUC
M+pTqfXa1rOyiYh78WvGjbAqDyJn83yXeMDG5nJ8+5ey/UQGBjTcAaISQPfoQ0DhlyHiM4AzH3nv
XN9XhXUSq+Q+9Rp2s/lDZGM/7I4Ku2uisG/A1M2cJATcbFZNKfrbH/62KOSV7NvoGDMYuy1dfUid
yq7vGLig9kAulMWLEGvVK2K+/kOfGfqe2BoWYW9202Hh+EseiEM2UDUwQhxIoQUQlrQR7lKT60Tf
/6vH5kzQNbLioupN7ZmCWjxiDdFM4Q2b9hM0ja9m3S+4luOq5kzLn+wwNb1P7G5Gr5RTTtuQvtKA
75V/9jgqKNlgT6Fw4SxIkWpGMvNs8MS7vwudhCMcmBpRsDZfM13p/hnqeU1jVE1A9OMLfQam4m6y
vUZ1M66Nc2foXUZCpIjlf/JDnEPJ4unjeS9pXbnC6dDulx1H43tkIgWA1Vp2ixuqpvMmucDQj9ot
sTODVUMMlNNUgLZjwVb7Q63BGjlCInybZzDE4LtKrDvM0aAPx6+ZXq5x5DpG8TR7iaTFUanzqJTZ
hni5DJJKfbyM87J9gN0U73R1X7D3JzoQPybEaQXEf6HDWDwj7yYxEbHTvEYmzg+N2Z0X5ZuBow84
DhN/hK2aqW7Orwzv1co1yfpPwIkzmM57MYcuhqod5uWdxvpN+cMjSAQlH/07qD6TMlh/PwaFK43+
dY70EBXzxhyRT42hFvfNnADSWnu1Lpkz3Y06cTXsYt5WA5BHznFAuAV60BiDv1co7hV3oK39WUHz
xefZM+wQ7Yw3NyBxD90rXWz4Zg2O0Xih+ktOFiPWKoaYQxjB0JS59LIa2Ng5InkJkzDAT4swBWhq
ARWcCGrE9vYWhlsX+az0v4ayTLSkttrwoLDGJRcEL4MciWHltKl6bTbiw6j20ZNHYeDA4f0GLGJI
VpF2dIrFJeK77U/V30R0RCYLJ0Sy1YUxcoMRbh8fV0EHpw/WjXayE7D9XCSM1uppRnQU4eVfX8rL
1C/yDGDh1Wy4WueiJUufhx6oUAVOFIaZP2I9KmjY90SrO9pCmgd9lxs+c3qH/srzfGvDJL0sSy07
E7bYT8AL4Q4MVVhoHUQX1D8oM0y62fy8qJAuwvreqRnUrCd0mCdy1dpWzh2TJLZgJAX/QI5CgpDX
rUzMjLxwZzKopiTuNJoQCncXIsMSnQC35OmCV7n6b2WAY7t3WVz0ynkzoIZC9rZSSJ7irTAHicYF
yBtMKPcFIjNDo+y+kGGqwHxxbumG8yLDKt5iIc1/bFnDdxBdHAHXp2tHrTF0k6Nni6EA8CHiRqr3
aO0gTIcapxxMmRneG4vRdT2FuCDL+Eke324am16d3ovx/ZtSHOFQAAm5akh9OKZyFnyAde8FaVdu
zdiM/LQwLLYdehjjoQ+OHeLAC92/RffYEdMePSVL03Ow0+1BLo6kGsKJotaJ0yEO32XSyuZd70kS
NgTlWLSszfccfB8+Dvjn5O1kC7vzr6JAb/LDNuOtwRrXyGK+1RxumxH1Z2OTWEyPAvkHM+zUloBh
PshQvkUTvxB5A/Mc2h/KBppQfBqwUEFmGGi4hI6j6tkTBxRuy6Ow05/rKfeU3YK+byNCf9gP868l
V8NLUScaczNszCaDCGAQ/jnu4Fe0QJipCyGrU5X71AIDU7S00SoXLMzv1tcPLq8oCiP6uMEfZQJ8
6DO30sU27pwVeNaX1VyEVfyQwk2I6xSD2Rctrp0k2CpdksYwomfOofsmrbscrFcASom2PAJ5jYSG
GOrToctpHUzpAax6rtm41PfFzxzWZxfxabDkr/XkGE//GK2OYoec56m5iYousGTb5peJywZ+Tlhs
UWocnry0i/O9ryUodi8lf6RyFeUXj9P62nfQX022Pwl74E9KBSA+DUgRUHmAtbKcklVfuoFu4GLc
vA7X62cRzSIn8lZst5WlmQaXZSYs4X4jkTU/Ya+3UQf+qvFb8KEW84qz+C79q8tn+hpTUYEhWhx2
UAOdQuuVHTwIBEx9c1AjWSjx+6VrEEOdpkBTrCxqfwMWGwIzqBXXM5XqBPe045B5sE54YycjhD9u
d4BnOgrCvqcYHO2NYQfQaL9/uWEc4QpsOVpCQNeH6Mpua9AkKekIHkPz10M2345tCyrCdDt+fmTZ
wR2eO/wFvL5h5tLPMQy+kWPFiYypkoiFnLMq6jR7hrd0FdPcoGdTpBVrWNW8azlMN4MSTutRYAvi
nRdA5U36dadYgRC5tzcfLacrwLbiU9XSKqk/4nuJUKTPTE65GcdcZIWMB1JKUU6eyQWuKFsqcLaT
41OLAZUcejvfXOZVMZALryn+kxFRqs2xyS80T2psXqxMCARO6rljDpa/NzeHb23nF+eaDT0gAiyE
vdw37hhqDreIDy78Q2AJnsu/lz3O6OTJjfbi3hBmwJZAp3H7M/i5SyiG8LW6upbtelAmZ9L6zLM4
zU6a7zwwfuo4lTgC8xwqnJTufIEfSF8MeeZvNdEtg17VdsQ5oc1CRPjzXXMuWNnzMBZOY77GJn0t
FpUzUX1WlLo/+LA6WAwzunNwjjcyAZez81meeepcv5LuY/4tN/0nYV6FL0PG+DPBwX90/hirv3BD
aD9+azG1f06A+UVV8SW0QtOWm5FbKG836/y8GobArPlSJlr5D2wNzXBD2SjpiqithWLv0AvWje4P
rMmZAqHJa7hIxNpwMtz9Bt68ieotTrQVc+6HQ1Pdnec7d6VKbHfBwQzr64ipQ/GGHjuxPx4eJp71
odyZTWmoQzg38sLAQacD7rZI1R8AimDLbsWrge8CubGQ/ROKS2n/469KZpITkfcutSzaDdSB4R3T
Pseo3X/jREh5uXeenAw+FJTdAI6pMcVFKL9D1LkpSCQ8MaOtmQ9LI5W1SVvnIQqdAEX4xgNlLEXr
rUqS1oIjasiloyi62gil3qgDxWEpdkFPnH3qST6hc1Qn8HxdYHuS/MQQH3SjXGCZjJXlOtoo7fdt
bf/JOvlueWFVxLwY9hojNzd6Gj54ykhp3zO/zI51KZ6RTr02RQTQktBSxgyy3gu0B5rugv7j5x3t
Op+fQKtGy2DiNR8m9zffPcNHfLVp42bFuv8GuYZQgYwO3TQB0b13DNrTE5ZlM0ku7FDk/Qcx2FBC
sQP5PRNYcjGTalF9LwhNfnq0QBguauJ+PNo1I73L9ih+gnZj/HlDuoytZOk9DcQtbZwnZ/0M95Ze
xSudkT70ls6WnjAdmq10fUlqjyOiL/sd6+1fbnREkV4OPSJnCNfbayiO49tFt/PekpTYA3Boucef
wwWizMK3TTiZA+JBb60GxoD5pVMVN93LH5ecIx46XyYEU80Yd7DdKabhyRRD3TH6ay77qM8IW7e5
q9E4nx1VnJAJj1OncplpZnin97W55dHBZLTbsO909/klS/ylWFBluDlguSwASFcryV0E/rWqwq5O
gQCTPKvvX2ubTywBSMtBVWizq5fcFRW2fx0gF1fu9teEp30jbJQ8M1BuV7Ld1Nd5nFYcObtBrfve
GlWFcnhYz4CiOfg393gXx59l63D3sDSixld3qW/+7NaUa5xS2xM/WBA9K3WOsblnAXZS49fNuZhP
O6oXoDwqZwgXIg6DJKGDIKUj2pCWM85sVV1d66RU1Tal2devtO8xTKMsENxaqL70xgYIb1wHYDxX
hP6tRqIzDBQw8HDMlDgv1UD1NkMbKsEnmnqkdNrHuxwX7TK4f+pxVzo/EdRI6rDv/FMcJHenZHc3
jQrcjCDa/EMtqCDbduO7n/KUveFZPh6CRIt1e5qVxFLwKbOV3vcJPwlgKyseTCIIShzA3tCazWLT
EDJhUKqB9yT6mqaIN+UWDmzw15mKdcwqzAKcH6S7NKe/GrFe32g4JiOTdi7R+UAdCjE9G+chht9L
1HQQYq9k9fDYcpXClznKVllhtQtO8PVmXEeAF7LYnQwQmpV55HE9QRb5ElqbQTfL90WQOAIpSW27
hB6pkg+oe0TEYRm/m/KpHH0ES1f985ufVFxn2LG37wrPnL2pazxwVch6+yRh9ZdawGsG94Z1BMAw
QRAu/TZAkVJKx0mwFIgFF2HXHVuYfeZ8Vw0owony1+DYcRJLKYR9INpEUua52YdOGsWu6s+KKwIW
jBTINZTMrTSPvu3udP3SdI4eOkdr3mhEyigiQnYn2yqhNyL9DGjHAUeLmtZYajEIyNpZPLMXVV43
Djw41g6+jHLVO8gHuRJbPv2CT9Fjrpn864p1EtfRuolQFJRh4vitHAxwryPAEc8Jd/qBQGpQUtaU
fEhiWPSjdeyxChexjaePjfuEnGiJXho8LPfcvilerUHQUi/IM4fS3yNn2GmLc4tPElY2c0fnsCn6
dgAT2PRftbsrcHvJlPV/5Pj5CtopD64RCisplV8OJ1K/xsHG/ALvT63+woK+ndO3dEQ8U6p+ceho
0cb3sx8bdj3PGGBYcHUM/A+Tl1yHGYNo8RP7ut1nQfX+n8flVLu95FBE5heI6ktmVBW09feaK6oG
KMpKpd746QsISj9Vz7PDhXTmr0gADu6N7/XU2ohwAJFwq5ydeI5wVyc5WXFG81MhM12aLbNFYe7Z
7w6QBIW+c9GBnG96aImXV6H8CNvOXzicNUU6qFCV/ri3Ik364iHBydZM/6ajFED5O3pYUxTeugON
NkgHO2BDbjYVXqH5qHj99kaNJhpa2sGxKz30lXENNrADrXEXgKBsNY9ZByA2JZhZhke3VBqsvikv
+qRScBizbwwM7uMNsHVhdgG4jCovhXWBIFUcP6hKVl0EHGPoeY77uusk3y97LSM1kW1y06fwVdo/
xmHwzKeDFG1XHUHIPVoyzTWct2r4KwfSEWcD03wqggCmAM2hDxTV7pgwMlVmHVbXodCsGyEGAGIU
bXi8t309TcmW1u8kHlXNj7UsGg3Re8M3z+0Vr0USsnnD54vZHip+0J9vYbbG1KYs8lOJKNVHAXIr
ebdgTEkC7kct16+saVwb1tUgd+8rLiPqelF+Hkk2F6qxdNoevEM/WbmOgPgX1f9qJwIn4g8MviJT
XzdwgIsxDgIR8PWSrquVCYZ6GUqityd3cQUZcsLqjmBTN+2D/BcIYWSMJdX5pe2oFTQFlNO9j6GQ
5cKnLUqONdBtabE5mrESppvzNaocsbe0FdnqmBj/dDW7UE+GuDYwYnWETPQcDme2EsJvMCsocuVA
imWkz7IlYAd2Y5I9yLbwOJBCyI4vjLdKGVwUJdK31VBb4rELAhllWX56dcZH0BgfivNwMqcHbdQw
To5APtT5qufmGchDEbPJKSkMwWxn46g2CSi4i+bWD23uFTy0ufJgtTFGGCQl71rgiDzdG9Had1SC
auVJEfUW+Iyy+XdPiEZv4cDK5jpP6Cv6OR37ELhTZzmK1H334WUdXvMHsAMS7j2o8qneJhF4XslO
d34xH7Vi6c/ImIiZYrGx/MyVUS/ZiDLJXgTC1eJw4L6ozkbVnPyZHUFzlIda8/L9XE+FxeqZfHl9
IZP3ZOgvzHmqViN9msthAqf0x+oqowS3vXQagQFXncBee85IYwr4p9qb50aP1JHPT002Jq/6bmDP
+yvm8luK2vx5TVTZ/ZfA106dil/wDYx2qTR72jTqZNgl1FAJp57BdQbyF4UbdCnrBuPkTOFiZv4C
93yo4mvTVPlVsdG2hR2BVU3hwY3RsBvXEWJ4OzCBGZxiChU5rTsgP/ueslTvD0Y0Lgkjet1q5bG7
0FJaF9Mc9m+TerIznv0qm0qdYcb6Wb+mQMWyZlga9rg5n/hc2sDHYqj3t17OEf5kTKOlUF7Tk5Pb
DmMTEOwwM3uaP1HRA8LWNKphA72YYCRj6WdlRhhNo7Y7oAasuyLdBSx9HztNU7FOfkizEs00ywTA
BC4DJ01XlxVyhFdzD14RF6iy3NbXnoUo5+NB8l+OZz7wv/x82+AMCvIQzbz9tmBOzSEFR29Z/+b9
j5BrIQj59hnOw7qcE56XWnvktGIWa/9pXNpE2h53Eg62Hgsed4TfSPIzEyXnH1TmfBb+bmDM7tHI
cCcjRgYDYPaIkHkg7ShojfSSAG3/hV2vMnH1s8YEQBJZ/G44Mr5arxthSCTg4d/sfK+3b1w8Wz+T
E81xSjpV3IBbAAW3U3lR5Ff9dgSEDk7xZ/YTN7nT0dHdNHRCiYJ3xqyx1q6qfgyEHpUa+V7BgxB1
m0RpXJUWEeA4BKn/jrv09JQsrSQClHICt88Ex8jV8Z/vpXEb0Q7hAnFRRD37DkGALQdH/luNWtV6
O9mxepUA6E2TApr0IWNmpdhbm9k1/iEeiTxc1JO/vNbixFMeMjEq0LLyDmf2IApuMKJ6b8PobOjZ
93Kpe0qGz5FeCXUNaPgxxas/f4S1m4hcc0aFKoryEDcERs+fy6+fiDIY6GYRysmLhPKPKdugnITP
Z2m1n61dwrukjjQXcJHZexgpjs+wNpFzPs6AckUzDlp/JJuq4Gcf8cEiqiUF3f9SHZrUI3cZpuit
ItLVwP4gZhL//FBu6tYSDdCAcBEkcNMal/kTZu2G2q6Cc38MjtpJLnQNg77gSKIx0Zg4Uc7RGdB7
2zOJoIzOifNd1Wk+OPjVpYg6sDz4YiJA4bG/jcJrkiGN8osIbdbmhMUc7YE0i5C2E0AC2UZiF6w0
uq+ZZyBzqz5V6NhO4AmynIs7NKgnXDnNm7/YfZ6WFXzw1ZKaSw1znlpm6k/1gjODbBzsMmRMS1KF
Rxi2pZij1ti1Gg2vOvcNgEjpPWjkBqXR787lsSfpKrIBtJH88gKHcZN05ez+cAMAPsqFelTc9PIp
MZTLM5wdVdyyY+fLMIzn7G6WZ3DCIkFkmjNmtdvu2UgbnuMN1S12W87kFrgPIXk2+25caUHAZQVo
VBOab1x4P83mmgOruIgozrsIBezcxDg8wNT5WDxVUcDsNqJvZOes5fIpQgIhTorKlhA6GBXIfyXO
QkOv7pwD57njdMx/im6MHxsgVvFYT4RA8JJBmPgt5qPSOUCs8RIgkJVX+FTIpj7yoi0+2snw/Vt2
2wwlTYtfm94qQ5/Lb0V5Ui14p6ejwK+hgUnSuF5a2VUMVtJb5Gtsdusb3/R+f+AKTfRugBZZ2m27
UNFf7Oifd9AQexqKiApCZkmp1uuJbHak4O6IgNhvWwChsU666tC+6ZhH+ys5tnnNVrXlHegkLkIi
nEDkD0+hAXniTH51sj+tmnamXgAL7EX5k68Fht5aTUizYhxjhGyByfY1WndGFx+NqrXxMz/qBCyK
PuBZfdyktHidc9pQcTkLV6uo3YLhwXRG6ERiP+hD7gKv3Wwhp7KKkHtx17LzbApw3bTfvpWaCEdR
xc+Fel9dO6QxRKFFVs1gkWZ26MaKeiYJhU+dV+xNhStWkF1amL/+vRyGjPHMvTNWqQdixTkXS0Tl
brDB8WK7KgBZu2UvShwxbUiMUt6vK7JXz0mjvSe68YtUCazHzInHp//esCHZLdqhNqjS8OATU1/A
UVfDwf1JAr4mQoDeAiBvbpBF2MpMlqo6TSZkCdjc3QhoMiZ7L3jkr9goYBX9czHCRzPXIrsVGyw4
gqQzFeV/UxdvW82andW4QeZmrOx3msT1su6Bn3ZV8+9aImAOc79FI1hmBGZJDZLsL0mf/iBqGTek
hg50E5291C3X0O/oPiqoXbqJSeG6lRqiSzOwjxMSkGy63jCtQEonNElPm41bguJeKQVpVI7726ER
r977rcqmNrRCCHl4O82Adnok+JvZ5hvLMxmfDoov1pnkY3QjJKN6Gx7S5MaZJpUrUQucMdPCTov0
qKl2EMpXpO09oKlnwdkslpsem3S6Gu3BsAlGKOTlGznVnhOC7PX6fZpzf1q09NNKOC4SSbPL4v6Q
L9MH5shWL98OaoV82E2hfttDDrWQVYj+wAmjbvDR2C22iGvfcl/Jp/bcH2soXJB9bTHGNJ0JR7mT
n9uTTh6+2QNcDpXiZWxe75rp8PqOHsiYlXxDxcIlKNdMQh5Ic7ZDGXDdEA+7cMmSOjamCl3TI90p
813my5RPd7xailBv91fFaL/gmkPIE7cDe7r3mLnjDS9o61OXiHqdhzSNjELqcEqjpEtmRQltw268
6EvzxoYazA+qt3GCjtZ18YWA1Sy4uhf4Zc3ohEpTnmTFrfH3q3SyZqHe+hzINwT/OHCW12xBPZRz
4gcUrMQ++JTmBkOfAAbP3wQcvt7RTWoR/4XYmKqQw/UNRka00W8RiZSVX5XNKFzTH8kURxJrgtfn
k5HKiPTPZASLpgnGrrv7rlCEjKasJnK0kugo+7dDCA70W5IrtK+aWDkj7G5Vwoj7FzY5K3o+KcAL
SRUej3SyH2LjUf2XvNS8K8dziBs2UGKdgGsg50RbbJTgElUT9GSuVfDXX0Y7bIRrKJh5muaZk39O
xQUl8Fthd7ux0mFAdh35AyJjXKF/3NiUh3+9BC+h6Gh3hayijYgdnKn68duwgWnPWouYMGgiH5rr
5hWryTSA4GWTF7996OxFuCjbXM47Jsvqm9H2/qHT7xUAaDaL/SQ3KiKobO6JtX39u4j2fE4/ostj
+Qc/rQgAkWrNXr9Cvch6tMIKZ4bIZ8UAla7vEgo7X3+Grtc9IXJ4FCMk0AegKK6FmpIHPOKQG/c+
TevBEgp0m4A+ZpO3pvhwc4mEszHMYfkzcjKagAXH2E61b0/kWXZXorrMx+R5mLFLfva1S6Zta8BW
KzrsxlmSGrk6WBgsZc033J0giJokvBGtvKKKMQisH/tcQ2H7Z/NFQQc0WY5TPtgh8OT++FaY68RG
8yH4OCvyedzf9s+EekqkyCSOgY6ennlL9Yi2cdfm9wVzn+puojuUpz3Th5IlFq2JA/Zu0SfKdxjW
DDGOuNZK70Qx8FitfnmwQe5evLg3jAKaf6+TNnYlJPvW/5CZmNatXbwTDoQv2WyHBAmWAXJzTXJ5
tO70S1n5DeFhjce1upcxgk4jbBkLaluXgAuns1AMTMrIifRy6mtxd0XOHyyMFvlLr1MSQ8SMNQsJ
lvmOjMAk7qd3gNsEKRuBPdPfglmoaqhAlBsSlc4f+TzO93SKq2cTR+3KX4kAxTFv2CHjLEnbaS86
TjWqyoJCOzgvYZqj4Nh2q/zYuap+k7b+N5WdhR1t0W11jdrsTY/B48cIKWF1DWjDVhgEBs9eponM
/AWQEwk08Ueku5FrAfAHLvxIEG9KRkjGiXgOl/WTiTRTd1abVbqukWSA8K2qH2sjZjGAKxUyZp36
phkWpPrGxHPnrzd513ILPJ3VBI0LUGB4BAOEeaeMVXSYciVlUkWu8nSbq3NttwJ0+iuY+bks5Yr4
iNil0yh7XgE+GDYc01fRgicGxW4I8r8pfKeRtjgxrhG/0R0psNds9V5r/WsVlx2hZllu7//AEg2z
Nn2Niw86nMt3euNljJ7VcJlGnhJX3YoE0UeAt3QUjOKkC18B3ZJGEjd0Ko55QkeGuzN8NSN3maTI
uuSTa1jpqsFpOhpaPmgy3JZH/+uCVGJ7LdZMJWBeswJ3cTKsM4RLYBqGOqI6TRIN6OSwaB71leO7
YCLv7eWM556UEwN1Y4hv+jgNZr81TcfgDX645a7M9ga04F8sLsttgQOem6G81aVGvpRsXf3L68ob
J9/IKm6wF6sURp9Cd4204/lU25ZzfvPGGakt2qJQ7VolWbtMFykjAEemTk0IJfAccslr9kZXBu5z
n/4NNNepGTF74S5oQ7O9wmK97nXs3GnZIUDL2aUczQswNjmhlRvcWsaV38FI3Iv0eJqxreuH1ujK
Ag00blXYinx8Pv6Mc9g7BuTJQJj08DF3fZqxscmHlkfgJfXuv1LCTAQKQkUpZiGksYyJ/XYVvUDv
xGkVPdzl70VEhIvBR0FdOwe+Njh1+iycGknPFBkRHSy86P2ROj0blBlSRZAkNfZEahVHRLTvbdeS
yCxoFvc1WVR948wAMB05YyXG5McCZdjfQ5gjcRFYtjuVk+dBZYFH3A9D+4XkJ4aU9q9sRtGdG3ba
0OmKBuL5dSzfmSORbGReB20qnYmPYeXu2UdQIuHH1Q098zOkej1KLOsiPyf+kuBoOQf4mFkJ5h4L
rO8SCoUseHS8G+OAw3p1RoeXV3Dr6wcqKB7CY2yjyaJ6bqVfxeqmvD/FlC+bN/jfNGAlvtJAe/iM
/c9lamNmqfHLXAh35iFNZQe7Pk3vjgm0a6V/PsEzTi+JD19V9TCqkfW1L0sciZ4Ccto+X/WQiROC
mpM4FkBwnZVZpUhDPWMVUpp6E/P5RPVyBYbMpbh1OLQek8GXoQmQCjVTw7WUdEasFIaTLz93l+ha
Y0D4g38TWfLJUac7666wLUpetrHtVMVeRopbED3t5/fyFPppJI2B520uByleeR0Zh+XynmgtuWcp
vC+ytZZ+OZf1jzi7BwuxCvAlWme+p16w5faCiQahJplVpsElgUVCYeXYBSmdtW/55dIdl5Y9Tgyc
TWb4SPE+XnkviTikXAiWX4G7/IolXD/NuhOPTNslqCniXe2yfCJEKYL0qUuXaFKefu0J6vGKmIB/
V/GoDIz9pq2nLdum59ewxe/Q/5WJFEOdvJjW/mRnJHm1+ZKvZkB/mpELnvpBwnQ5bJaoABoR87GM
N/tsUlyRhmzg5s3emX+ronXu53P1Wdirzay8aQawhKC3sB5D2jaUqky32HtTozUDeIt7hAmQA0MR
eFzAlkxp7mmioUkKMNbl8JgwYVP7skR4+v1BxSQ1yWa4dPOjZqyrZk5mJfsvDAvCYlQSV0irW1e/
ikYSgZ47KJqInG6kdAyOpb1v32exadiR2E9K/DgXlm4RQ+Zi0IIsiEmwYdV8p5JwhSADEPWLkyRf
zFrPwI4qxRX/mLOt750HiaPfl8hjBXL0NUGlylGJhUQ8+JwoIFtCg1t3EJ4V5lqNXFUpy2uQteSz
kMqUwapXPiLY8/kgwvnqshyHliAJsfoTvff+7H5PnLDBRUP2Ah+M9fovgG1THU+FFo3qi4FWToSK
Ph85GQoQb/4dz4Cl5tc0K0bSvsE6RgZrY0BIYjeivGlrcy+Kz7cDuV7fOZTEB8c1X6t8RskLTBuF
Dg+H3011XHG1IwgvyDw3X92SMIOi+1n5oUHpSkMa+rXMDX21cPd/vnrgWhEunV+sLrwO6m1skujF
wIyUtvzJBKOAgs1hvLG9A0AEGrlPuz6Wiuhud/pMWNO+ExjmD29yyxPbS1h9v1gNKZX48/UeXh2a
qyLDtb78dn+5b2XWDbx3tE5aRHp87Fh1pTK6lF6vusLrx3uP3Kgq4JwLfwGio+Id1nDinZPLZfBs
p4gLS2F/ZjW2LAJhPtgzb0D/FpGdPcfavvcvfcRdrS/n4PCzrP5irGgf/plAO5dZ+ys4N0FcmJ1z
pqSxaXqhUQrb4u+gsmYL8pVA0Gf5L5POIJvs5IAPGIrAbV8h/ZuABZ99s0hIHfCWl2y8IFx/CZ/+
0BKrvJFGoQdgG+u2ynoRN8I1FsJgy3epRXL191W+oz2jJ40ZKcw+TwPHCmv8xyArOZCvagjzi63/
Q61lIn2Zmm6rbfvVoIMmX8Aa+s/2B044edYx3Av2rwR0lUioEs7PDFTG8UF2ePQFk13eBbxh+vfj
uf/I/dCSrCnY+dmPNWcgFRQJACmNZ4ccMBgyerIleWWQf93hXhVzP/5FgYXtfXvpsraS6qM9rYUv
hFYea4jCkPwoLq7TFNLuPypT0F5w2vFyfEV/T8777nRWMl9uXqE1JiF+yXkxLBgkb2AnXu/378N7
p6XpCK9n9uLwDKk66SZJLJIJC2VmaWCG0Iwj5H9qf66N84MXm2t99Mt70lVCq/Gv5n8BdksJJWR0
nqK6ppld5KoGhBipd3VwVcz3hEM1WGYARjK7Rw0HMdTQevBvM2yU4lX5A/4vrvBNsMIw2OO9/Gun
en6OKUtxhU7uXgN7k49MjNtSaAoAzigTPEVeRP7B++2M4q6HwGkKTTwAugiMXA5Yc59cz5SelliG
y0TbYsgTKCbsYh0kOAjOSARm4IgslDFTMzD79sllFuN/BR+yl4dDRJ4DXqjFeAV/uuGxGbiPXU/C
AJ75t/K8mKOFYvdGFdElxpQG0iW5ih/zSdEX0w1s9c6fedMNlUsoafqHjBInIktrynWK5YcmrlY/
ClSZdgoV1vPI2Qk6hNVpwYcZubf/jdf4PDw3uP5NNWz388fdK4an5hiNwjoMJeeywRD1Ki1EGe6e
ZAnEO6+pdoDjL+4WRvdgIJoDHMILG6ZqkJ1YklBQPciPQklgUZ+kzovRXietnX/72GOacRU8oh8D
R5BTHskBDqG3yAumIrxnPGvgEpvLnA4PRJBy4eb1atZnysgpy0ltQEjSJWpwMuNBCay9aoJiFjek
/PnWkdEnGv4vcVpfvUs6gzrCqxCjf8xn7i3g/qhPB22v8EL8FlgdIMkaxCWKcHtl8gUKHZz9oqTL
tW7irXkmuXV75uO9egcohsQu2lNSibY4BS8fPd7LgG3ToKUtHPfNYz7e4AlDUeEvl0pjUsYlQfaM
j5XiMYOgeu85b8kTlsojzql4VRvhnuhwhYNZq8t6aLjTS5MQTdZnvEjo9BWQ+bPE0Exhzie5YqYq
It9COd3cFg9Hwy5hVYEzmrj+43VcucfZVtKdgWgSAAZkAmSHhXqU3xfaLfVZL1VbLNyw9rvlCvm3
VJfZCapMtwN6A/CTHkyxz4uttGy0FQJrMWWgFcA6n/VrWtoSND6PypOlWGnqwZ9tfglEImtj/Mr8
L2VV57ba/RXmUjo2ij+Hoou06YQTp1UukpPG+Iclry0E1zmUdMgdCi1jMbme+jnwRT3Qx+re41qH
0KJP02kXXwa9S6hpjRiZszgh14a4GD8sNpvW+mQjuaUCAnoMaJQ3Q66r5ZrCZICVMPLLcH84hlNb
2nsNMPeTsaOkZVPM1GYNJ49Qnws+cdYnhNmOy2EFHCFIEMwiCXDMwYslZPNJolPd+b1Ejur78DRm
d480QfJd2ROULbOLdOhyDvLt6TZ20V1jL/2lZwtBEZ5VnQT9eIYhDFh3ZaJaQsVqNJPjJAyOfai0
qy5ivM4YynzM/wZfnzK7hHB/8DhiJPxLby5W43oAVbsGF32MfRNgFU+Dw1rtoemP069R8d01O6Vq
rcV9itdhAqZ26uGplVKhtuhiF7jK5KOQDJ8dH35fm2uk8szLFIdrir2LOVBn7tt1v4+9svAUeXHt
vcgKDvfI0pfk6SzLzAsNIy43KtcQ8rY1yYN2JpPE4ECOrh76Am2SqtFD6YSFJbKcFv33KF/Nf4d/
JhWFJPRIyYNjxv0gpd4oZPwzzpBILTg5Z1myv4tTZwvH6IEOlDj6F/bH5lqb1jBAfzh2Ltyk3j9q
5La8BxqekUK1NlM0z+S63lG6VMqibOD2cHDjJKeN1T251JrziqbGPulbos13W5JLqPfJagZaquti
JRtWePv3i2EQ8a4ho7DErEYfoJg/htXWlI8UIxv2YfJgzfB4uIZfMyr0WbhnseFZApF4lqu/LVCz
AX4HI6AXYqbD/A6c5tjzdcBRqW38+3QLXo0AJchS0L7E5kC/ULbrPC6SzysOFCw31Fmjl0Qa3PfE
ouTGg+hQwXo613uL9D3f+x6TQcQBp7sPYye30V2O/HlPcErZeJJwbU4hpUxF2ZTE4zn3JQ0i1dwJ
ChuBVgoh2Q3FWEdoHeOuab9AnWs+ZPl75hCxfc14b+YJfRTPbFXRqRT6og0FcINtDP97pfufublt
JWscBhFU5YYQDBJrtnGA4m+mZBOGMTnEghA1uClbds03dmn4Pf5JMUS5VsfvQD5MKyqOt/R8L2Hp
aowX1NRU3RQuJjpQo6mpjdKEITwNwtSoEnk9pxaB1OtSha0d64fXQFEGMMeYJPb6+25OBs2hjdRe
q3duQrsObpywpPVjrQKvsKy44j075HflwGpzjkOXUp+/gwziY5vLQ69lu0KKcGxUwp4xY2wHfdo9
g/q6jd4kVHXRtB10qyV05ZHlE6ngR79OReCHF6A73m0Z+tSuB9DSoA1cio1dv5w9I9RK4OOX79dY
HlqBFZZ/LPLPnzjbGMFdUzQcb3ZEQ9VGyY1rPJsQu8gdUzeYWYCbtnwXhdr9T1o/JZ6CZVm49vrD
w9Te9vNPkrU2u1qrroM6l5xpSNLNIK7955W9qziMeCsWst8wBsaz4nkUuGMsQXktdXr02ji8fE9A
MdZOwFVbkUhGEv7Y5UkEsehhOT+9ahrmh2SgvxkeqaPWG6cYnLe9O8Zrj1h1cOoSm6EGns5lUe8B
5Woz5hEk0FXiEe77xXOI5BAi4rYHkRYKELTOAJs9kogCGTDC/MnrIPOzyYzLVgbpc3krWNxbmSKD
ldDoWXN9GUASaN+G57Z2sFowkHVr9eA3bO2xPc4h9N/pnlUKClpFHohNv55qpLpGa3nwwIfkPeSz
dlpvLVbdXr8gKtFf8UGoX9F2lK/zHgwmpir/7t/S1k1fonWJIGv3L969O9qMZcEiEABYBdV2w4aW
ScUEgX8Q8Aevx/Uuc5dZnCoETvjASDDIzF+YsVQJRrlJOKNIc3BgX3s7e9V5/3i2vGWEop6SAOtK
mk1e3HdaeCIRX+3wx3kgSWgxO9nHZl7NA/d9mwfh8BE/Rk9lWjpw60upW2yodQ+XfqgToTZpO0Y0
xevdt7Lp5pKQruSjfIcEEyyqQcaf/NV51i5ptkMD/ZapSPkiBENLHSmNfSJHAuro/NxKY8axvgAb
NzG3HRxOWV7YSSF7GpkRitrVHXwgcnGONF+9FZ/oMaAkiqAOTd6PB3SnNxzAamPOHkr+OaJ/OXK/
hLL20GN4qaEI53F98z5nnrC0QEkQtqNkfhaAAh615IzGk1+gxm1+FBx/eCq3C8Ol0a1atgdHVySO
gS5VonY40eI7uU1PgXMEazo+N6Z4FMhpHLTMoW+6n59+yF+Atf0+0W8mhZak8rIR2DWsvoItuUOe
XaLvpKXYCW8HcP36OO9Q8rBtrdR+9QL1BRKPehxsZ+stXFUgGaay5mzYsBYhGNHQCNQZWJTiDMp/
CochP0ogH8bnDPijxME8HqTnXfYvpe59icEAENDZmXtd+C2HVNWIUB7bf/Ht4rOF546YGSikaRfG
USVJ2DnWSBN/p6Hs3FxtmUot/KGUrlSoKRNhfGsNaRHgTxF/MCGahWya7VzksgUH1LGLblV1J2qG
urERHlBqZA3ybaaEhChNJjAh81MX5F41xHj1l8Bh0qVLtNJHU1fEqu040RIcV43hECwAzDLxnUgo
l5isIhfH117j3KimrPqGE1RuMGPyOZTCalEqVTIE4g6lBMRC7eSI19FT8KZrliHJ1XM0Ix1JJktg
AuBTONF1wqIv2qQfWTO3yxDBAzDp6cNp1ln++SyFsGomJKDM+JBVXl6m9AFLtEmV3NCWC7z5elzj
6YN1GwqqnNRsU1yaYUFEfdQu1imT86Ftqj//xgMo6OVVKpUmIO4VAM4vx/b8N2QySjcco3d78RwH
+3jyX1cJh0hyBkMw7qcDkYOlawirR2w0ZitX9XfY5dr8GVxV84u4IsA/v6jkb5rSHxh79bgLVC1Q
ffU3F1YDL/FZ4y9FaEomEji7lX4FyS9RigJ7doAIK7cQgTtA4kYrqWxBHwABKqIb4eCMZRTY7b0J
KkZ2bV18v1XHQ9FxPJt7YbxmghxFhN2Z0lQyZAeHXogj+enpWJymCeZWEAPaEumnicVEXpSl2R/I
rLpQ3xGKbHWpVeqeyoBatMsEusmQkBHk3rth3V4g0iqAOvh/BkmgCoPCru6fbADddzKEJUpxmcpL
U5dzZoqalkMBuE3Xi78j6ZzYQfQac8p3GFdbxx5XyTskfgikPf0iugOFfRJtg50YpLSAhyCSFDah
tjz6VjGKWAUNHhILoZHl/7BExy+SzbeCId+aEeUyEGdZTV0krOX6bW3UIIMonpisCjlP2hDhKcNS
DG7uf3N/6yxtLjhIiTa4lQUyoeiV9IDkcrDWPEhUqms3z7ENlnSbVWIlJackAyIqZcxfJq9Qg0B5
zZ4UDkka3haHoPj6jiLu4Ci/DXkR/dDIeTfPS8e7CysaCnHNbzYyBa2GYuYTUbqJuRJAQzt9I8hB
5vjqeWCwkWgXXq+/ZuMXe1gfeZBiObs7/ukpFBxz/yu2cro31LUz48gE55i+9GSFmGNy92K5bgx4
F+h6kaYPAlUrQC2HGI4Lyst3Zgau2JI0moymQQp5LhjGzH7zzfa+3Uhy1Kw8hst3iGMqGCnNEJkJ
9Nbm211A03N6ZaDwkWCjgeER6Zw+GBFdhZxj1xSG1n8yYThWiOPC7hOIadq/SOQQ1NEAXSPPgwe1
pGw2Ex1h+eA8+W9jwK0IGHX7JPoEqqPMhDXULssPpZvJ8kr4ndGWSQm4HrgQezPaPo7grtObRQAO
F8yforQsMqYBlccBdCjdcCu3FQaHLL25jeOiq7B68cvIxzG4yQU7S1q2c5bZCUWLOo2x1taF/pa2
YQIgS+1DL6+GmrFdHI/xeh21s060MryqM+6bA0Ao3RGzpB7axKl6l6BUjc1Kuhj0Mej83WCDwfj1
QGgwOEQgH631wvLkGPHhoefJZtqyIovJ4vqyszb1nPpffNpKPR3TwifN3el8ltiINIhghrqAlyi+
PJ2ZQLEIgolj2RQgfGL+rYJw6Y7ayinvGeWr+UfQ951BBUcEDsJVgEkdCMFvVnxujCIlVOgV4d44
KnxcBXYtXuvayOCEAcm0f1aeJ46NgtC9yk8LlZ6ZrqMGIunv9GNLNz18ulQLmmqmAQpSgk/SaWFL
4IO41+qFIPKDe2VnHwPIAJFkHwNQ8p5v7OH2+6B1SHJPn2HdWZcuOYuZnVRPKKpHT5hVOi9BzhTj
3rLnrpkySBk9+GoszRRJRbwoAiPJk+dTdWmukcY7XxzUaxjghH8SfcLEllNrYR4Qajan8XlIqX+D
r8n2LClweU1rgFz+JYWYFSjF5mkRD8Krq4E8CFZsnRdK6ITPH1USGG8Pe9dx7CGWWrJtkGM/DQbv
089rAb4jq9N5PGx8mIa2m8NEaVRHhGz00oPXWxcev17zTwQr9KRcxK4c/PypchhQDE7a6b0LQZPY
cUnC7/qVPwK//EJYAvAfsVvct37DfZyzwkcCkJ32IDjzefMOl/iSQ/bedb/VW54q/Jy3JknUfJBA
9WZYHQljm6CPgqTN/MrgHsVxb08akbDrtTOdr1ogIJTwskH3XbitMVWei35yx2qvxGFrHUfudcAy
Kr3+CTFOE4W0CmduHYkYrpZK3Xk2yflN51AT0mz3p84qp+xLgpCGrw4pr4UL2ekXNhJgLNTRdMxe
j4kRX1OUAG3UzzaNxNX5ybOTnCK5K7+OHB/WohB68lV7kiHLht0ha5GsC0/WFaH6xKe09oRrNTKs
DIrj7Xhiv+ES4/PlINs4ZG52wDNoJvP3OpQ74VhIfJY0LZkAWerM4afEPRxh2ZvbIbjh/IO0gs/+
K52gd7XmFBQuFE5aUuGgYy+rIklDLOr2e1cWaB/NAN1Sc2iFrhLe6jOCThToWlzXWtgzailZUqYK
A+5pgE58sL6MmFTk7v9cKx2Rnhgy2H+GY8nBLHgNjvJqAr/uOmPnpWKdtMvdwsSChYEUBijBJ8Yt
474catFwcXTDKNt1ND4KE760x4NlNAISMJeSSddv+coeMovZHZ/PSTPcSXBFo55JNSsl8lvBK/gm
Fl7Sdkxtf56zHcZuuMf7aPXl+m0Ydm2v3tQfB+MVSA3+8NlHM9u533WYihd7Ii4KhBgzN/zHrUTZ
n5f4j7L6ePX/8jjZhxibNvKYeUrJpznsQ23vC+geMxiC5qE0YARk/b9y873FqhtyKqnM0LQNMyJV
TfqdVHhlkrNf6JbMz57EB2ONtETPWFsq60EeiqvAHod7bt8TIuWbadKjWQ/pFsgpT/Da/LQunBjS
Mh1HpN30rCrAWOp0fnwHLPDXuCULBRQCdFLqWe+Cld6LL5JkRhxDctErFEigDlkEWiTftvfe8zWy
gJte74bX0tx28Mvq6DEt2ZJTnjm9H3DnAe1QsJCR2oyUelsx/chQx6a0pd2fuMdDINoS1rji7eaq
Q7AwhkufhNHa6GB4opnxRqxLAF5+MW0HFaYTApe5/N+S4Ea3zZtjvdB0q9klNRouV5dfGcZo29ij
T3M7vbkE2GC/mwyRmgsRIdSvLbJEpybfcz455xeTLFecM8ZHvhvhqV64+7nxv+naLY3RL4ebqy/w
IEjeDbF2cKG9+U51/c6X6fI73VQzT2IwqcJFpSz/N6BmkCVf7deDbsQfqLN363ydd2s9ait5/Ixh
NPMuIVbxeMElMYMTu5VGewCdSEFi65DBBY+Xw/nLZaCWqggjO0H+y9QW9/Wyrw9fl4XWh8s7LIhE
5yuuo/2L7IWcrD38NtutImLGwi+0QVJI3RXPSRXEImVqbbtf1vPvHJkWGM+hhj9RpQXArFjuCGpm
4mPHt5+vi3QqY1kDEFBVffo8h/btTwXFpX4zcRacSCuyqd/Phd0aJQHrzgAFfOsDtz0UWAq1RYJs
yA2/8PQCRyeeCKcA/BRUm3hcnC/6wlagPicskeFrD8W1KxsQfJUTdRqGVImoscc8TaUWEMu20dKr
LPtFaCKdH/n6e6ZiJ/lIdRqDG7nA4JYIFI7V4mQ4PuwDTfCnUpVn3nEAzq3qP25CJJr/SNvfIXWe
DK+YnXM+JQSoRecUqyZjY3iW2K/zfUn1+c9CvJSEi3soxhPb1D1qZW5VXB1s+AnJMYeGY3GwNzeY
P3wDiKXcvhBfjjJ67bg9cumoycneP/cg5Yie4l13Bh/LPZQoANkfn2J9MXhabKuJdiPGEuMEY+Uz
ed4fZwxRxgYzgU6ssRzbi1S5PYpQSaKZ2oKpLI6fFbgugC1qSAFTqjoLCRGJqM5/ozukxrU2Tf27
Y13p5AR8c4V8TohjHDYen5PnPZBZ7bRMrTWkdeyjlSB2e4Ou0NbcYikBPrlHzySeBOveeCa13sOM
2gxvsF38TKYbfTB1WX6tDrxwsz6txwXDkX5QJT5FKI3L7iVV59zV3PXDocwdhiWeaR/XtlWqpThB
gFtBtUl2EGK7PM0oZy1ZB/yRxEkao87YSyHJV6+sVAYVumLwH1u6Mh3puL0axTTyeKB/v/sQh2x3
Mb6vSaJX4fUpB3C8N5mVzq+QktirJNTOjRrDSZIDT22NVZTo5WuIWM+sgUZHN8257Crz0Z6OkBFb
ryh8ZgQ7pLWTINoSyi8a6A9DwQKqwKmAuBiK7PX1wCm30GlxMSBUqFKHC159b/4Mb4c5nNGbLQew
8yWRk5rS3kkd15++RDJ3Hz7qQeKN9NpxNI82jxChpSKIkgW0X3giCjuaEcm2AotdGuVYdxc8d5Xl
TM5INR9WEKDKF+x6VuGlYwxGJp40XEY0HGKdiWv/jLqeLSAHmVDpiMDwDo2BldYa9MMLq7fLBo8I
WV8AdmG1wNzTU0PKYrrXmYkOB5NHXptMR976nRE1oNVIENcdhVWBYvs6Z1wznKmXo5D4SyQxrPmj
ss3s6kEFeEAwgU6ucgWSHiDsoM9sZR6sGh+rV3n8j+GfU8LsbNMPcMnitoGXpr3kvaKvpf3YxA0s
NsHaQfXRO3OeQlCw5bpAi1CjXQ3LAmX4qlkOAU4xGBRYj0zkdbLNH50EPqJhLLulBeGya/XT7Udo
UVxEKt3Ha1m7nlx2PRkEham+1lKyeOxvP4Bnqzx1ySJ9N9yvlmbyGdrpR3qK3BQkXzsWUA5LfGTR
miR0QB4MGaXYMlxgJS/i+B0LMhdH0F4tjqXNBRENd7ihMvKZItyRFn4pmYgMZLXW4Dna4JakrDui
Y6CdVk8dZyXv5f5nIlWprwakEJDad8tRChiOWlP7cA4/mDAA78Jvg7pGm37qZnfIquSPZF0+28Nz
1pzDw/C0MSQCGZ0tAEaUMlMnWm96Pw9fZ3KT7g1aXbD9FqzuV/9Hh4YM44uWa7LMIV49OY6uzYKq
L7qlAQ/IfP+mnZ3oWkWoSadEZCRH6b5S2Hme/LWTBAhjbL0EkXes6d8V9+tOSRYMob7WfUfg3NHZ
INGNY2bQQtPcXJJW2IOO0zA9ZYs87i7aLRyjeoHV8kwx5eTLWeZH5/K2ngZjkaJi/+1stkesbZE7
7jz4YTmeYZwJ8CKSZINE9okQELDefZrbrG6wsi5yiR8loEHFRO0vXLbL4UiCad0QSgp/Vr0bikeD
IV2X+Pdw5M8t4fcLI0nVT6BOgV1hEbPxqVDG/Srh6qUfA8KZKy1IWpKXtZZnOpx8VzO/vJGXg46I
PoOFwQiVacddXmpsdX2Ktgnlx5agTA9j4p0XUaIDfuZFSXXdbLxWAgyVBPLbgitQV5tCS/wo3XNf
/HolRMnLzfaJAP0HhrgDb89tPxrZK5qhnajgvOrfVAZYGwX6bXjTbtQO+MMyAXO0d0lKtUFTv/Ls
hM6OnynP8OfCfS6sCgjk3BUnYCpqM7xgRzGSKblCvgyY7ZA8UnoNSmaPkxDBMhv2Rxe6rTj/xf9M
dnSWvSFI14eDl0ibShONwZWT0o333xdHuZfVCU6ov1FqAUMUF5jUd5B4DkDYnH8hw5Rh4Wgb3Da0
NWOcCv98AVs1V8O4XB1pUgVpVNcUyvKbmSA2BZHaZyKDjMWfPQpyS7YhCdgkEz0YiwvdSbO2r38a
v5I4CQilS0vrY74YQlfF5lQGOlMDQ1S1Dx5KJiWJUotQlm7wLs3eJUEq2p3sensFWSJP76LAGOFK
rr0Vv7DT5eCxd2Ge0uUo7Alzvj1Akx5lriV40iJ6ydZj/SF+WPsMebACMP5LucWaD0bjB6SnDhkk
SdEFZAPBLDq1wunxCyKAlahBcDSE+68l4dOY4NXWmmJSDsPjUR1auj/rnVaOKOg8hLvklb2kZBIc
0fkuTLjXvNyrrfdmvfs7iHbDKbVdeDlyldzuL5l2KBfmrQ1URCDrWgRQepRvlb4gLgro3unz9hGe
vx7aKLmcXZxA1l75FeepCpPz8x1SKlwfzlQtPMVLd9vIAVk06Ejhjx2Y+x9IHMulFBWY6MaLcPpu
dzB5luH1mql8RQ7mSFOTjYw1YAOy6AxQaFC+zrRgeI0D0yVC5b08utIXVJE6OioOILaS4jkJKMYM
mYsLU+1wlBsJYkgKZY4m6MK061SRSkYuCyiD3VhmgcGALMVcDhsk+55Mv10GSXBYxJ/2FxBaK9Mv
p/JZkR/OmVg1O9XOhvtOyScXnDOMiL1J5oMxSxsBVcgCA/Hc0ST+CbUXdFTQIrVV5OuIPlhKBNqW
InjTguCFzlbPZeoEsUm4MVp2EFnFbO4/uonvPpIAokx9vgphuFpzha9oYxR5dqo+kkt/s3qokcdy
j460wOo51rddO2YPPeZwKWEsdD/wweSY5nAzpdTMfwWKM/yGA2Zak3NpGgsPdergnDMJoZrkOj+E
Pvc3PaigAF3WNGsGOqttR9NvTtitzfEpE08b6FpRhJSCgky4K6B9xI0z7cfl+3O6UoD0YtpP/6+J
X8ocWCOFEfHA+4LCHBT7mR6O8I4ahWkPvE9MZUO4Yc1QelLr7x1GFmIoUhfWvq9lzLHu03pM7j5l
ulRt2Zx3/coWY8atBeWqk6RVq93CbxLhqpdyIuN/RhNgx0PFEihgB7oetOhYsPEbujQUYHMQIB4i
QZkTKQwe+I4G0vnGvQ42za+0JNZBmVbTH/NEHxpT1MfhG34ocD7puoc0f1/nf8E4isWSuUk1S1Vg
v5S99TYyYupC3PoqQ4lnnmCJj/nyNP3Tip2P/S8IOxZyMcB1I3zyqU4YBxySdR3r2o/TyenacSms
Zh4X5L1zfbSWBgpRgnv2EyrMOGn2gt8TqddUGzOTr/lEAL0vWxfZek07TJNjAE7xjAC18wS/GEK6
YkKxrnlGwPOj+dj2aDYQBY+dvKzoFZT7mK1hkzwyeQFpj1JvqXB6d/pmVhOEpBEQH/g5w8lJX9xD
9p1p6YGSEitzP0gC5vxNgdanNkj6JfwBzn8e14nD9GlvcgVq5RhXbPVUhtrsClLG0UfF0QWSXM+Z
htZ4bHrWqXeUhIqKaeH1jMjSd7E1tozb1U4F+AW2wGS/PYVoVGZh42sD5qA5dENBNU3d/ik2lcJZ
L5XdQnvVSS5IDVz4/mtqGxSjfxX/TgAaKY6SqTBi3MiwubkIO//EQpMSqsspfAquKQPrIW+rer5B
+1gY3KFEYUV3WxWXJ6JCJE7uV2aiPyDxtGq9wJUAjEAH+kh1Y5p81dekAh8OGlDMPnUWhtdqrE4f
9OKqNheciMFywOKpnVnmarDLniWrHP4qPGWMdL7NJG44ov3DBgMOcjlvPcohj0ivvP/g23QfKDMb
oeikybbAi+w9WJpmq/X4MYBY2J0/SZ1z0QeUhdYt8kaxamxxwBNK8z5pl6Q5jlWRk7nr8Y/r0T3p
EUjHs85kkx6G5QaTvD0x/gG4pd+9Nkf6jSeH3auOlZtL5Md23O0Bz54KgxIXl+IQ3NhRDqvSKEFa
tUORLWYCi8I/sEr64XxGp/s9tQME2gFm3mFSzgFR6QFIp/lJDr3z3eDWn8psGmgiY83ewducSjji
HtAUU1lxX7PQrdN+bhKTrLuuPAfSgm7bef5O7DSD2SNYNCtitJLuFbeNS7aukJgpnbMSZFV3FccD
Sd+DsOtrX7faHT5G7Wwy81rbreIR9J+lZO1Jf0HMRwNeqshyAo5fDP5D68kltaL7yJyoRp+tiAaG
cxGhk22stiy+zQriNA4jSL8hDkZfRMpS5oaHnM0SUJeN/0OLrncevfwwbHnpiEht24Z+yI2DjzVM
8mdc28UdxXv5c0pdXdcmXvWpiKC1zSDrzRSEOq5wACnvDQ0QuxnZSLZ91gh8ENHlULo//zrVPhRc
7ntjI4FnS6dAD/oq7/6DgXHPFmrWJ33BrblA5/sZCSt6YFdqXlJgbiJ41iRylSku0I7t8eaDEIme
qzalUbhPIBCRKaPPG7uZH/6z8LR2sxOa0z3vkHaVDaNKgftLtnz8wrkmvu01A8NLN+/JEdNYIt70
+9LWtn5mBsWb2RPbzeoyly9a5rXjMDp+/hQBp4LRso+FXy5QbhFae5FCVpMV0ZnYS7AeYMs9cwFc
AGulf1y9SUK3/VCU1hkm3PAoYY4ot4A81M6K+Yshx51b0ZWY1CZbh39HNOfphSUWOY6yI3xl/UjC
g6XPKcePpaYgjiQYoHwYoeAYNe1cJMjiAxtiJOBiLqF9K39TfNoDl4YpOxqBEWu5B3ovrNTc8loy
V3upK3GMpBt0GqAZT5lWIpJB1pkHvqZOq0l9isxa/EqqiZyJwPh2lCQS/ecKbhSsLYTk08hLglkx
2nrQXTFdgG8cOsJrEZgrgVxplNMhNsS2eq2l2uBaii5U26FocCDRc5hhvmN0uWI1Uhkv0c3RMDiJ
npZ/9xOdHwcRvI7BEFT/rcSRycyaRl0opcw8iubJc4+8y5vjMY8bLZv6D0Qw4FZVEPvYVo7cJdXQ
e8S33/jPuEvn7Wa0946EPzaaxas3W4qxpveXsr13xSSWdhTBQH0IhEwsyom2TH0lUpOYal7c+n4H
D1KJp+0goqRomnP3WqPaZ8oLkoUO5+qd24e2/P4X6QBgvllzmwOT0+aOZF3ckUlLaID5qH0+d01z
z0eWwt05YIJMIM8auCnH3Zx+Czaw5ZkmxqQEIIFUsrtYhFjjy1Lt6SqBib7/53RS1BCdjvMQTuCL
66gg9RbngivW2sWpMGs1hvmpcqfEXEO6bEys3Feip4Kx5DFa1et6bXmCA03oyQrjs0Vyq7MFJgkE
iZRRydU49qeXamYzjosFWl8cwht89V6xKh+tRwys9aae1sv+eVKGxhoypNB68Upc4bRXlwVMpxrE
obBVg7UUnf5ClTH91MxWFXqSI17tVGg5amlMO6QrDmuaDfs+ra/5m/bYqLIS2XiEgCnBN+BqWgiy
w5Xbf0lCPhhkKUx+0QawkioPQJLqRhaVzI5dEjQypmEsvWLmGrr6g7cXOjFdHSEch0WhVwCXCYct
QdrOjoTf57/ZtraqDEy5ddBegRURsnzYTDoo42un9ZyuocWtXYBz2/X/m74XZzG2zPa4nAUI33sz
7F634oJRhLhOk0NSxkJ8oSrkG47T/eEvZ8vngGoZ+0vjWLnEyYyTaRRQUDgXZoce85e2EUM9TJYc
OQqoSihNTGoESALBDYPaiU3aGZhXuZw+krdZPX6tnzGHPLulor8YoudNvvrE5VL5jxs5RwnEgd7M
ENKHKB3x65H+EJ1eiJ8Wk/11PcZ80lTONQkmN0CJKWC1Jep1eRbYf9N4Hqm6c1ANK4f5ovGcC44P
ivfSAuf4ROXtwHoNnlx3mYdkRs1www6wLN1ImpbGqaEndiGEZjRpIfsM4qUgWY2VlQoLJ3SFpd+P
i8dUXZWJbr8JrMcnUfzniUPF5BvX2FX18E1IZo49tD4QCBmg5SBQ56k/wD6/Uo/XADouKBrXlnjv
SHsXx/EWJB+mfQHGBs314Cvr/8PWD9oszP9Ph67nHivTGXSv39bgMVFHhHPy7V3r4BkXetEnRhHE
lBM/gikBzj2o+hhZzwTNPcXZHcYGi+liGucrFGSu36nf3aYJDk/B+9ozcQWLIQNrISgmckm4ZSfX
MwCIvagnNgpLGjj+RGqM9TMhsNU1h6MNv9FEfaMUQgA93bVidjfrhBo69WRMozOio/Y+xRQ2/QJ6
1Z53WaQWwJk7Ls4sth6cmpwdxrVjj2Dx4ae+cpGYyyeYC5BZHm8XKAYSXgDe9IN4CXmK2TMo92vA
PpG37d9u3a+KXc7KQZMsGoAKdUUhjHWxJo//7Gqf63s4zLlLBhBCmSU0ZWmlCkbOMr+Ak2y6ffld
7okuG9OuXAj7JX/zw1r/chQNf1Ix6xun3nE2wBsEe28TnSUvnNDNQAf5N6I1gufESZKG46efqSeJ
nZogswyjAtotngRMfYi0qm7HfpYR7lKA3b826t5gDRiuU3ccM4yK64xO6rWMc83VipdlzkMsB9n2
OSJUYICjNfpTR1nWsdjPpR6eGorfAfRZpDiffhaViJx2g8P7gvMWaW/Evx/6ocV+Mqt2pzMzK7Ty
lNC15kDA+7YO+27kvCWTbo6q9NY8C6mvZS4faUCfMo/qjNYyTIFmtjw14nOz5qMWAkRr7qKS9Ukt
nN/Ihbe8qSmKzhM6WgfE+Jjuyf/cP4cTILUluiIkAjDyDmVsZ0gkAGrMUX3zUU96EEN6fCvw8NkA
YfRMHPZ339sW7RiXvZMpuGPjocnad0ccPFnNhIkm7rgta0mWiezQ8h/A6vO/GxWKbmLiXn3ZGfol
F9BZGX8P85U9WEWfDgZpSOOF6BOUuiEJKW0zruzkPudedxh78G3UVKf9vk9UGi0GGBalALJDfSPx
hMA5KvLw0Ws5ivkIPjHQHFLyYpxVnz1Ru82jgE1pKv88Z1/Xlo3kjRx0zcgDHPVeQ8Nv171DTyqI
Yc/EfBUEP1jufa5OPTpjt8rymj6fmn5yhfvh/yG7RoJJsTF5y3zRVv5hCgzwmdecleT4u4uZaS3v
8vb+m30WBLzXxRh5mHeVwWuVDSMWuzdDScnZlXgPOVGHp88a4iq1Y5Uh0LZ675MICTXtoaWbZhl0
X0px8Xjza9tsUBrRsyytlZOBdZ95jyyAhWEGkRW0ma0Z5KNjUnLztk5Y1ja16eB2S70dypuEFU+M
//j4b2uXdSjkgP4HCIqsZSFepHwMI+g46R2SIKBlkH9zAIZf3d2SD2yTCr+HOpjVCCppTmqEH271
LFZoOdPjxtPLqqL5XJS6khG6HUFwvRuCe2yrN97VISh8DMk7fQR6KVnsCrIpWU1sJj6xtwHKUv12
YDv7OigGgxvpM6bg/SqRHGvcvADy14I6F8ENnhwRKCRBJyMOVNVdU7M14LfxkXEKMWtw8/mkcYbP
rnem4IB5tLuiwmKAslMiqDuNCinKbpa1YW14yRcZZRYi/NBruvYN7xsQ8a187v2EfIuis5MMNVIn
VMAwZgXW1kOA39Ntl28YI0WDGqQJ5ZGi55dw4tSF3yospywcYMq8q1HshLz8xDzEFDAB5Yfsdw0n
Z5dVVJXgB/LSMqSvKO389Doe6i7/EZqTqJG9pplxISGSFCVPtcBsyvRGz2ZZ0LMczLYM2LNjmuE/
sO+m5XwNWcrRgsvLMJfSjyJ84RfnK6E+VHONmOquxfQMqO+DphWYJkKHEjATvO3S5lR6kgB/XkQg
ed8kMGCzjBXAwqkQDeI7aucHj4nbwkwpN/T4t6SEom9Uzsmn55u9JiT7/hekn+EF5PIwadfaGRYT
kTMY1dtUksRiD02gea4uXY1lknydu6wgLLDfYTQR9SWPSxQ7HIHAP0KZtnAU1KXPwnZRLXVbmlKQ
ACiR5qbw4ciTIkKr/n1b1brVFlA8GjcFijGFMHG4yH36pP60p6YXpjqIHrqZ4ZrsMnxNPqPaIPZv
6PRJ9rO9vxsjiMEwo2YDCKDDOzs09widMbNc8jCfyzMe1H3vE1NM3lC8ccBVl1cEMGH/PfIRPtDC
SyqVHgZWm9FxV1I5eeriPPNay6mjBYGuz+8kCpOJM5Qk88e7zSokMzXEATNkjqSZ3FNjHhClRDGc
gnE1HTYE5yuzz3Trrhvzegm/mjtn+TeiXmjYxTcyS1VnWLgW8aMIquTZ+96fuBt69jqr+zbWXiwO
1M71/q42GSEryuE21aI9nUOi6LKG7ZLgGf9lMUbIw6e9rYOKbYFitneH28DWkBcQytgt5vK9cAyc
hdb2szyQ/lcEuYBBV4LfXcBwopenBow6Jc+MSHMzBvLuuPSkKSG4XhrR8Gvdz72sXEneeU8yFXj6
IAkjE3SxwRxtjf7SUzjBnNE4m1iu/LvPdrvswJ8URHxwAsUn+63HTRbVm2Lw0ZNZVhKIQTTBAjfD
7uLm5r6nf4r8f/r+fJYT8O2mIpwbSNTXzhSDBc+oSKxLrB35zeb4IbhU8chgs7XeIXYxWZ3lKVe5
c0UzFHcGLKY1muPlhQ+q7/nUrCivQuYCSwlerV17zmiTNQFnxHtDj/68aT0Pd1p4E+sultEnviZA
Ycshp6rB32pg83ctgyvLjYPZ2qTDJJ0K4z1esGUjEAU5eYzfhb9458+WHWl8XBMAztfpgs0uMkVH
6j5nWTi/VSywzzGZsIma55AB8K60RkSR0Xb7Nf/nC++hnrM++MyIyqhYmsD8V9geF3xVv1+Ob6nc
otXlVZb+cVdp1P2qBF17PkZ5t7CiAHMgYP602cFIzAXMys78+lus/pmx1lIE0cAD5+VO3l0c9hHk
WxSU7RZQGOIhJgGfiygDgz4dzayEMZE3yQppa17VJQDhD3pAoyQrcsbTlB8vfq0VqxhN1yEaWRtd
MpC43jUGKh+q9863ZwY5zETY3JUbsRhfS405bC6kxz9LNja5Y4S9QxdTWhRpMgIuU67cu20IO3oh
K+ilcJY2M4qKAMZAROJSCNPsxWuxfE8MpWSjCb1fh8JQVqfYrjXyz2lB9DmfXkCgxbe0pkCsdNb2
LXRFG4AfcqfgXmJO5brsUvESkMYxfBiy4YdK3/4rM70vPu8I2xZp7THpDPR3nmSjDlV8kRcSvGPo
MQnFG9IfdiVbucaU6AAeJfTeaUNjxNtFDqPB9hf6IcLG4mT0CZExFQj3gwOf3BCO1jialhK4IOTG
xuAYUXxM4ezgkJBvKwvy0nFk19WvEe04au+0mIR6eciIoc2zcLmPF/wzvq+d8JIWREA7Qm4yn0QB
0wEEbSSiqVA22m0ZXRSsDc/k2ZHkR3z4dINX+ySKv8Pk0WWPOeXBju/1KS8nM5SoiwqP1rIyVhS0
BwH3hkIQDNV3SairXzwPByM8vcxPd/YWHNBJe+XUguqzuHkFB6/6dmRlMLqU02cxCECV2i69lDn9
bG/2OS0GoMp144zpTPUX/7dbSMO8EkiaeFTBFFocZO353TWDAfaMsjH8sBLB+Z07IorcFsC/KxW6
ks29MK3i9z6HU6caNJZhh62ujxdow5X3S2ch6QGAqSJhJypmVL1ZxwAoqOnLJ+MxzmPki2DO3Mu+
NpnuX9tUqx+JzWeONDEIZsMHm53ww3EFlNhXAupVCXdCTi0PYmGHdblY+eUpGYSHwLQkhdOUGFIb
Nlos8Wr7KtdLR+8HJMg0/DnPBcTam2DMZq7+/YpfI/1P5Pt/cH3hmBYZBEdavaiG3DAaGZVsge4E
TsaJ504YSTeogxehU5d9mvfll27XrLOvoDX2z2jgaOSTNqoIOzcEDs2a8OuFB/1ZyJZgYACZLR02
REs+vqSRgmd+tJ064lU5yMbLhlxBjl5giB6idL7Oyln5foQ/5VlrrT264gaSbwX5MkFo4OoWm0JO
uCAckXj7bdrs0UdR63EslnRa5yRTRBZ/K7SQ4nsZt2DRbgaoaPBgzDB9FWUwMtdqbQICJBF2EIuV
Fljwn3k8WRPD6ta8finjxjQ8AI2TfuFjoO9BYUphzfsoKxzZ9Hf8y0nFk8XHli0kXeaOhgdxGE5W
kwK1ZxuFj1gIhVkq6bsm2OQtTVZfgKXMs5r0w0ZWpiV4natM1UPMp/qmN30l9XJo66aTFiMVNx51
u9spHBMwnuGQDYs9+CAbNbePaOSdGO6MXU0D7HlCKoQRWx9MTMZ4NbeZwkHONg5xqpUHss9WcPge
uF1hwBMwEaMZgXO9OT2gj+gd8RRnCikErH4TMbdvyiNnV6lMRPl2VdclZGDKC70aqyd//GQRgBdQ
c9sosNOahbNK4kVEjwxzxzahSuTiwe8FGyBTAodXA9tSfq3zTQ26mAccZmzkLjEkAnwhbO7TLkmO
PdevSRwnWzokqY7SdW5Okt3sj/J26hHhzvSwC3uw7Dq8e62YT/baZSPkPHvSlZnkdDTu3gVU/zvv
xGGCvXDSWEwqZFfBcjzwSew22TyZYV639TE7yJ9P7bE4nSADDkq5co2w0Uuqto3Jg8U+HoqbhcdC
iBely6rk5VYHUWmDs66Yp1EaqEVxLeUnF3DIgcrJN86IUB3Mtrt8dqkeuSqDMM1d7melbsZzxpk7
MpVYoHSwMMdI6h+s3MBVr21OFBhdIyiAjWQG03SyX/JrkOtldPgE4SiBhGFgwxk6C7pXSC6qwHC/
aDomVgBPCKKo3wqNQbCGAOTzSn51wE8rGFDfK7/r93U3P+cYjt1eok/bhW9ckW3uYsf0wrQiToCF
f9WVQB/cgdNLMp0fwLAuDay0rvpMDO7BPVmO6l6P9YwTlTBZPXPb3pgecuXypvvQGbzz3o8BPU06
ct4FwHHXhWUdTQ65adL72sTFz8NuhFYnlfpXrB/mmn95MpDGx7FTUWknm9JhP06K1bbgJ5A1JVkv
lncB0RbaGdbO5DJNongezDpRS9qGG/22O1+ArxZNapPoZE7cFZelpRZMY2KiwZYIpWiJFTYZHBxI
jXIxv5pENr0B0h1WkSOx6mShtLfP57vjYKoCjxF+a+ffYpM5Q+UBOieDuAlqR43one9aLV4oWwws
AsYiYn1Vg/iYJG1K+2T5gydMArRYK6q5WRK8mdCj+EyqAPChrdFor3VB8EGVqVbqudvrDJPeteay
+tdeX5mW1CHxbPUiAoLJnvh6H6UzIoS3ahzK7kUFqAWx439Qf2j3dkJ/8Qb7agA29rR+9Ellbobf
dNsURc8wZHpbRV3R1CKkuXyUBtK80Tw1ZhwNs0UmVRYh1t7T+s7hbRbyM6AXvEqvF2eT8GVxZByT
CO9Q/RSaFI0QqCcG4p+eRr7cLf6KvGqYpTq5ZtU7vRjFoJFcjx0pQ/Afpuiwngr0XsAG1y89YOtE
Ds0Egz644pV8ALuXCTHFv4SEVas5ccx8lxo4FZjUgnQZ0N+n3ej3/KYeQIYZz5OW012XvUGNIsM6
C2489mnYxfnSPH4xiwhxmUDwgX2oFluZnumQ7lLJPKGnmqfxG0jEOQBF57YMmM8O/8EfDEOcVKiV
lEeqv13LEkBbDm8AahU/vDhCIo796WRud41ThjQGn254izBF35iFSKPpkaDgMykhDdUn5DiQmCKL
ByHoJVPGAOICbM+G8A/fGZG/FGby4ux3V4BB4FcTZ1alOD3PLlBIosSYjob8QmeoTzwwz1x5I3Ek
ERMjL0+/Ws+nIXBw9L/T4XHDPcWtCf+Km2GTpyBO3/j2PIBWaqiAzpTNnuzWoBOEsR3OG2z/sFvR
ony9hNka35PfGWYYklCWV2gYSVUxYzyWTOTUIB7sL1vmz2Aq3RRi67UMZkAZ55jDBr/k6mHgZ1wd
QqWrS55O1nQ5hMI59LRoViLkUAfs3viv7KHIhqwnPi1bVJ20WjK2AFfl+Wq4HMEtPu//gUlexroK
mdGILV2MO5XVQO60G28ERWmnDcMCDoNybojKeichAQHOR1SwoFuj4ExUor17dMZVV6cg5wpmrvCE
wsijNVizKPeXgeBatr3JNLbT6Rg2UPcSTw9WF2fuPdUKcFSfAhd7qfYkbNoqid1JIO0G2ZhE7Yxn
QeTrAx2HdereJW3X7LlBalSeDddOwKukc5ielUOehDkJibcF/87wtRdsue2IGW/EzOM8se0uf5of
btnGShH1iSjzIeS+WRFBafO+FVn3o+xf5F+OHQqk2TpzBmCOXZp93EhsjFXyt9q+CXnPajgpq5r7
mtinS9GOirLqgK5oySGVnj56ewWrpz7hCpKhzTkUAjruK1GWBRAv8Iz2lTXrU6YQE9w9Zw/S+xBq
VhrEyBrH+1CkuOJOACSigeI6bjddC56cSsprstWT08po+SpEMlQWpEfN/WR0RzejiG9NwxuNlTQS
TV93KXmOIqyjboUvy+syoASBm4HQ1XS+ATwaIDHic7R5yzz+pqlO7kNqQi2A9aiHS34vYEz8kjBt
wU+3R/vpGBBJc/JlagsDa5P8lOGIcPXM/rdBRBp5I6nF0yKIOgeoQFRn7dIEFJ42lgywmk7tIl/s
RbJuGPUWX+lApGafrXgFeeDdX6XscwtpjanQrYaykOUn/FI2Et/CXtcUlijSk4R238rG11nxY6YO
LEZyw35ONkgzjV3InfgC35waOwvinnCcjOTeRhnvxHrkHqgKyYRW/86LFiQItLHtA5OKevzuEM/d
5g1eHXS0++JUt4OkhShu5DE5+lOvAmabQ0fhGTqBy9okyngAmitSnwQMxViAJ7NuHL/ernEqr/9X
Cj++yf7GjB0DDr92rXNKmheP7MH0l8pkXOTZGdn1YEsiNH6eX0hl+hzi/9MWthJgCRpaL6aV6SdK
s2rZfXIKaE5Z+DNn7MuicZkxmvmkkZy4MR8wZXXHaGT+TO3Unt45lyPKbY+mzgaZC/2BPr4vdhT6
twbrCzWn0Ry+2jY4GfINBNjwt4Dq3t3e2AXBL9zX7Xc0t1+RC5oRDXLzne29taWraRNP2oq/pxaF
xyM1N+7xUFZgKn+5S9tIOWJp+bRE8D8ptvRsejTcaRYBPKCLNGX9SY/QhjTqcfcagLW0bGyoAGHY
FnIQ0IpjsyhBNkZpJthy6ByyFDhG6I2ZQFiUopzrfUyPjQk/+EKmwhy96msrxUaYf4MhX2Sjsl8b
thndAzYum11zai1wXOqHBK5r91cls4vk2Ik2H7m5BjGajRzmjBX9wG+gL4bhV5Lo71xiC6JhUkwP
BeZqfmod7bzb5ZwOyMvQfq1hc1fd1apIGzFwbm7hBpARlUsKK4PqwEPx42YeAL2LvzbObUMRsWz6
odiNEeifvOrHqBfEeecmOKvINJL72bRQMj6JgsmZc87j2gToAfhO2IW9d8V1FFqnYB8t/9RKnpOh
5iIFSYsoKzKzm+nIulBj030Fz/tRvOoP4HJCrmh7Tmv36f0np6H48bsMibSlk/MKpn5FrYx/qGwH
3zfOPW4UnjBBBzyf2ew2TYR1SwWVfWx8lSK9qoFPRYZSITR5oOtiA+nlmFA4oQPAfBwYgiPIfrRi
ILlQMRvAMNaXaBQkM5z1QfxfIWn+cbW4eb6OYq+lzWF3OgzYMAsCzmS7Cd97CYmnPRacjjHV5wY+
VjYdCK9SjqI3A4MaBPkSKJP0UpG9rGMGM0Tu4wcetemcREf0tfUcZmgHX9Sbpxt8K+IyYqp3d10S
ppXVfaMdzaNWUl9rIzY0gc1zwq8LCSvCOnGQ8eb6Wl6LEVsm2IiLAt2GwT1kOPvhvGDNj6nEBCmu
x5IX0RtNAjUJcYengzj5oxHQAXwHllJ3z9JbNzBEZNEP6VQUKwrR7IBhANrycyV4/6aGYhOr3pIj
15h2+LjjiARKUT0uLfdM8PgZb3BX3xBl4zRdt10I7pgKGIKI6q/tGxcKXuMdhcvFkd0CgS0RhlaQ
M6s9mFczY1eC3KHn3rEBF508jj6TiRsIERSFZ3OOppNWcznQ1QBxqK+27YLqk+eF+8TwGZdzOX8t
goBcKTw6TmuJw8W5Wi7HgAWFVjPtG/Cu6xHTOJ6TFLEUY16Sm1wrdAckZGNRifTLFgZIvOJQMNSa
xWT8+HClB88toLxmWdfAuGt9p/jWbAH4MBT8ucNljYrtnrkFV7E1eGIP/OcuoOvxUk4LARSkmTL7
jLR+Zg/lmLecRQk8T48qe0SJYO37+xoVrkVLEivAbMkv47J4u7UGWVT5Jzf5yx3zUPYXHU4RCnoK
1iPofrB4OKCWkWNQAXSCEGTtAWrE167MNci2rquIAeklslwZQ4ZsskxCEwRycVfnDUO+AXtvhv0Q
t1dAHTaN80H0HQ7hMj/NXRKMxQCuxhMVb2I0Fey1cAxa/3BoNIh/edhee/vOBP8R3bJ6pTqSDuUa
sXBTkF7RCwX3IK8IQNt7b1rtBrPBUs56KrAbK63qFNowogXeAx9yPkIymqCbJZN7BIcjjlcm6eu/
y2HGBX2x7vLT+RqwJy1mLr1Ue2i34A53+SfEe1yAyJbA+nx5LZ9a4TQtQZXul6TGcQdhQl39DMT+
w17judE2odMjrBgHyeOCgvFf5x3f7cByJaC8Wsgt3sQc+sqXmhpDJh2sg4SY135u3tulhmUAGm0I
sBrPYL4YPIkFRihVmACZB64je7F794tm8CEsGxWLy/rGJ8/t+zhFt9VbU3YuB4f2eHkJMQd7E+n0
oA39a9763aPuJeIkqlVeyby2KTzPA0GTtxdyykIwF3OZHp9JkVh/k0ZxLtX0hzih+Jy8Mjf7XE86
ssAsPmaA3cq8PscwNC/J9D3ffRH+IYT/341GavSV6pRqRqX5l6dNfh1Ry+mfh0SIJTgKBpLblcLb
10kSKS1DZjf27h+JOJVNusUwzzZSfhfJ3RdWbgpLB7KhSiDm0vAaITSx/ju1ZZ53n5hOZ2hucMW9
qr4f84ln/7js0iBOuodG7BEwv2ZnDN5Vgsg01NhkJiiJ3NwNebD3mtV4ueQICb3ALUPMfYaT/Ipy
7nnjCR4Z4hoQDB+r1y2qbBqu5I5o1UPwoMHjNHoze0gASlKURLae9q2n9VCZYNY5dyd2zznBPMwg
b0qbRzK9OuVb9ZVeVtseOwAxCYdn7n0kSdRAd+fpf2+DBEBlp6M8QRmzV14HVJBSE9jDmPBDJXgE
sXLF3qyPt6+07ywCSOjXWUZer4y0ZhWqof4XYh9W0DJUcSCzc4fEYfFtqI8Rp7lQ7D7E6mTA/F31
3unPeMFKjkXcL3fSqxfsZIFP7gEBSkBdTwfxATjpWmQtSpH3YXLslRyvrorBwvJcs8M8C76IL0PT
cbTU50jNS/qvqdCgLYTvIW2qdatv9Zi64mdytS14iLvfc68LvGeFjB/KZCYzUKcysLaKwOKATvqF
v/cwosofT8fOgqK9zxWEjCmNRJZH7Izmm5mBT9Ye10sDDP4+p2s3Ez0iWVbVGSGaefUTYT9/ye2b
Dtfrv1GNimeQ1582TzaBRZIcrXGgYdgXxb5jbcN1WW1OsK1LPRuGbV0MAn/7evIVjM+Hc/HAcKn1
iEINWCwtN4BlocIJUCsmFD35R5IWnIxp3TWDrO3j07BeV6TNOcAs9bURRGC7PgZDfjm/GNiAs4RH
pH72hTF0LvWPW2ycvEEnlgmAiF/CTRXSZAEFIOzYWTfUy4yFl0vagaaFs4FdRalyWHe/vouF4joP
yYk/neJ9ol/hgHMZoTtKzNeoAoawLOeof/fO0+2k5x40BsqE2P5+m1o1SaGIHDzjYyyQ4srPrdRt
bpqNIiElHpq9cVH0i8pzqlG76yek1ClS4Omixvd5s5q0xiTPRq8f/PVSs6oex68G15q2VQiWkz1q
Uw58Ms09NbC9O2L+Lu83OLbyxoR0DHaKQ+hxH/mHZp33A0Usjb5oRdbl722jacorC+kpJaLf3ZRv
eieOMeVZ1gW2rSEOGa1o45mJhlHuYjnzGvdCQwWQEKyiNzkj/yaUE0cLqot3x6yXC8R00lFPxLFG
eWKZzBW2Gru1bbAfqYU9/vRrxkLbNT4zxYhYP+vN1YmSlEzCwG/26IIKtqXcsaBuiN8V2kx9TfDa
mhkuReRlqt++LRUmWd1f0oOXLzMbOjlpXH3iyPXlQ7sBECp0QF5tOwaWUfy9AYHEFaWqDo+XJw+V
bCpUNObqyATnkoZhm79S3qW2KlCCn2zEQyg7VAQ1tOlzjEH7JhFzv74QupXXaeagCPSFgIJQPjJ1
1Gnfm5qrazXmVuqixo0imTs3ov4ItJLIZ/erk4KJmeNYXR0lAve+0ZhT2zayjvucfwMnivsfw7jZ
O1e23eFH46BETGIwwUspTQ79BiF5vxUB316Qyjfac/IJ7HSQO5n7PkacuchszMTB9AQQKFxFw0xZ
q18+EABKJdaa7n0nOoMEYrLBD9XBut3aKCASY7/RSVov6VLE4rHX2coXwHE9CKuUuZXYdqlomOUk
2ww01HAWIJXpQ8yvFz1p/IT1XuGAi7Pmq5MkBp97pv/mC9J9PZVnz6O/blUc2Ya28/li929x2gX4
VTIYntdthhZ+xl9vX4ZPCr7/Qg3OODasevubZzTP5kyA8++dLnr/f3neIPJQrTFsAl8zWnXABG+Y
ddA7ZyutYDeqw+hAt8W7mClgv+4gGGHdX9Q0o+oVLPk2PTXJ/fWmXGo1/I4Cwzw/otBYvFGMLd7y
VndNa9z0jrzPG34oDmSndsNgksuYkrzBcGOmK5PbhAcW5bDE1QfgP30gg2yNNulqHGKxtviF/7jf
zR+Obuolahe17uJlLKhxtP64HuZfIDVAgxgYNjVv91pXEvZPBIgv4EudgYC/OQx4i+6HSqfo/pPz
N9PzlniJAhudOXu+AN+SqrKOmoOMDxauzVbYfnZDMLwBpsK9DEjmH0g5IoTTIm7vY2QY0KelVulH
IPQc15SSPVd91DxCRICqYwycIbIWjerKbnKqe1XhVP1G54hCBMGAfKrx0DXtiQ+f7A/iMnykkYsa
cQqhcCyL6iUgu9eI2dMz55thVIS8xsjaewxcPxJKnWJmGL8I8NZayh7dN/N7sMwJ5G+Cvn4cL1lW
IG1KmbV5aEhGaL2d2wtvyaxisovKfXvd+DKcXCk+s29KjTS6uYipNh2BQTkSmNrj/LfMY0FsB9bz
BczfvGYUwkRVGfbLBg3bOiO62/49Lm34nxjR3FmzwvSbq88442opV0LPWq6IzMZmp9iRYgVo+BuA
zIxa+B/4VgGpuuV0PRCI3J3iYwUfue+A2+oRtFlImAc93SH+yE6qSRX2Q3CKQomloFS5Oel+oZ6n
Pu1du5kSv+MiKvPt6NWSUWm3QMrz80EW8GtLbdeDO/hEmhsBxnfnBvDLNsUcof2NReXUy3L9kp4X
9AJBFNB1InrwUnOAKl5oilMuVtOzl1Ge9queIwD+hvBRKCE9iHN5/bHAsscuSjm7yhiqPAyeFjcq
01we/H0ruu7XMbz5q73mNSGNDC0NpeuhBNMiwn2VwxBEcYn0lzOjCaX5ICihUANRLkCMupBvKr0W
y7EB6gzXQyVJOIT3NAZuo2qdVLc3P/KTxgrI3cyJdXHcwccqwpDIDtXnL+fuSVZ9owq02p/sonXP
uTnJiVAPJPgEIf33L0Y6M9W7vg1+SRmg0gXwAJLLaDWAT8secBFBiu2aJQ2YULCp55u/oeS3p2tL
xdAz4wz0GDBS0jA6IkgEC/R5Uft0/Vfx51HE3+SkyLDO21E5AaBWmH+qxEzz54LudqPOhwyYG6D3
YWyMJDhSGSffnabhAmvkxEqwjsMuBsLXRRe3RMtlLzEU4xKWDOAlO6DVPi3LXQNDvMgRM1JAZyPD
pWu2bOCWIv20l0TsS4f2kw16cpEVTUUYthOlRAbRA5+mKuaMhAxLDs0+9e3mMOjCAPLjqQJTFj++
ThKNj6AauMLH9CkvUoEcAV3V14bnwUCIKtuF1vzV12roB26B6M3UdNAoLXSEAp9HG+5qfJap3Ue0
ehbbbBJ7D72XoSUFloEswBYanp+kAtVvfQgWvmmJ7M1p7hwXthNnLiumJyA4v3Hf6IP+gdRR0e/Q
sHjxvaLNQjqtEOHZPhDJN2fWyfFG+EdVqoGxZbjqXpsX7UVUw7/J46QKX/IEe0oomPCl1q0rcvti
iDuR3rHdWyOok7DpJD7gRWvMr/7xGoJtoc1anLGsdSaV4+6rOA1jIR9qwZ+DPgR4secuVooJsnN0
SZ41wdhqTF9v9fTJWfS9+SpW4FH0SYlKy6LMH+Ws6ZQihKvzX9oRtrKkn1AdJkx07O+CodmgWtoO
w6qQ/FVQ8GXHIV5ujKK0nOG5ObVX9ZF0p1S7yr3dkKC6TxPa3Bh6SY+Uwrmuh77UnkZa+7oy3XC2
62gJ2c1Cg7plYFxOzDsR/cP35Szh2v8Un9bFK6+/ACVxAm+kijkMSEBW89Q1Fkm4BzkXRL4TspeI
8TYm4HRLMFhE/7wyn9e6Q4MKQjBT3KkN8xayp8yIe+FNbdPZYez/IUXaO72ONavt26T10BHEtCFw
fuLdXRe2lR2hQ5CU+VU5Kcr+lrC8pmBKZCN+ZGEozHmd00Ti+T2QhVVB1vRp/QuuNW5nMIVnvH9t
1hKzlkLrheHz1JyF/BA03VzFlTBbph3w8f/XviabgFVDeHJem1eMwPqKyQTAQJlq71jmNsGQTTMF
W2zNeWO3S84t7yegN852Y1xbTanSF8OjQhSHVXNYQ6Dbw73Iug4S58jnE1MWCQUKsydNBT/oSipi
WUUMbCUYx5BYFzqrINKNBWGvaHU+p84hc/N63iFD7jgU2bXRfMidB+D0t5STBOcwKmCbGENqR0J3
4wXFEP8OPYzIa9f07Bus45XkGFVKK6ANwUVeX/ywa9M/f3dpW6wIupH2OEuTaKUE3+4yu3b9RQM3
eSE6t7EAorC+vqNmWOCBpQCh1Q70W2e3J+wdkjNANmaqNWbJqKR9xWMEKutt4IzaIBtjvGGtLu2s
ih1KRklZxiTFXPZDvvdqxpdwxiFAIJqZB2RS2ntPLDwEpYep4UU453jjDJaRLXVG9IkpI+OWs58g
Ee9/S/dwAwvNImUj4j7Yo4mcCfNNx6d6yPHDsha3Kw2Z0iESP8d4shBjeefITjMEWBEusPVgar9L
0RGFHoPTk/BONoJBmvCWkIC89vym9QpsyQ92yqmZhL8zYYLbczU9YwbhNp96UqYqkwoWqPJlFG7M
OFm0BlHkT3rVHj64kMdeztJnqaQAGxCu9Yha8amscJF3VamE1D/b1CEz4qVyN6BOycuLlBYZ7IU/
Id2EqSf1kN930uH9Pyxt6pxdLUS1jHjsRZylw0cAbi4JKxlIwwqLUvXolyB4TsVwOYWnDBbaSnGo
+NKE91xCfNVyFsyEIs+I0KXps/0pJjcymqfEO+gGz5Wt8oB0OzSu5F01UUWDcdRRkyZMIYommPw8
O/xpTfbNB0rCm2aE7OS0pVFiA/KTb83kXTAikbtwgY0ZIY0i+IkH8zZZq5stuKlSk5INTiUUZjdY
KUg3O31ZG1WJuFacv6CSaVnLvbEaq0Wp74d0uqRUagOjgwLfdYEKZA+rNRLlErdlINZGu1DNDIK0
SS4Yz7c835H45+uO2Vt5MzQ0K30qUT+peFLojHC8cyz3WG4r71KU8RsgZ9v5oWznDRC/kpOlhwcy
FERmpYb+zLEC+hs8q5eor73I80jf1ct1tfUKRkRQG/8CgyLH1eeMP+/Ij29W59Y6OBZOuqEI+v2z
DH/P0w3VqfA/P0AcMEgZjOFJ8+FRDwN69n5CFPHNCb5S2LKKxvEATBF8vcD950pQcLsk2QfmHL8V
ApOagLW7b6VVAaKC7Wb5df33kcLDXloX9ETY0UJVMhT0KvG9EDw+4fgC8Wflno/UpjfbXb7EFNUp
N5m7xm2OusAkq4eetdRViNreLUer2K61rXybePcePdQ8T0qjEhGCvgmXNVFxXaRcbkboZDIqQw8M
qzcIumr3nOIITweif0xI/R+xo/Q5awWUvPrpSC4OT2TYUNef7Kl6/MXH6m3Udcm9oOQDsg4M1mv6
V9T5WdDTj7AwKlCwj+AgJP01hsZzKOQ7LkyKQ5fTfFqSB821Qc/NewvcpdGmf2snkVoI7cH/uHOh
MFjwE7xC+umEk2AmuIsZy7HGJ3pGnzEqEUmSclJu7q2nAsyjqlIpeLnVD/2HKfK13IChp0w82YiU
cYsqfYWHdSlrfPFUww4kLdilIUFg19iYRW5wnMOI3xZARk9KaC/KZ38cwqBGkVlNzuQSVIDKtFtm
ptK3/a2QpdDWf6gTbdp3aUvZ3StG2+uR07SJgHdbAF+jM14kwSmKt3SW36/++uDcpwfmE8oqT8eS
+OK8RpndmaVkrzNagtiGG83FVZq6EXGQgc5HVc1DtpjkpjwqTUlCRUZFybI+eNTkbcxl6KU9sYNF
uZdHmmyTjCef/eeruLKHnPXdINxIvv0WqCOQMYjN2wpheWa7zn8M4XgP0409GhMXGeOCavA+YxQO
1KxtWvAzyj8TegvoMRpJeGc5jEC0Hiz+EgGbJfjlG5aUc82CZQRR7rki7SoepRrG6mzUHJvg2tvi
eyq9Kwlt7YX6YAliCut+vMjf4/+l9fNTrhLQksNr0xBJXjSibMu1aMfYPw528Nfn3ZIEmJcLhmPn
rnESPZ5n1Jj5KnFgdSctz9fAqTPlo3mgJQLzKGhHXjX5616YPPphZxA8DS3uJjYBzYfqj8BsY4GO
rGB5aq3Lm6BwW3rz7BltpWfJzvK16Y1ZaqcOGvmpJQqyHLXoY2XlnzeeX89HYlrTvJmC3eAS/W8G
e/RvnPcR6UM044NXE8CgvcQlStpj0LoMoGZEU8Uk6WcPE/ZV5qesOYkK2/9mLK/16gj94ngR3se5
c4eXk01zyK/i4csFWWmG4xMdJAuSTwpDsoG9ZzfqilUP+zdLB0dvXqJND6y+/YEkIgVYo31JTWSv
f2uBahueDDB29/vtt7Wqtt73GqdNQbKCxjE19lLdm4LfW+/SOrhBxT6ZPZNDGpz9vFbOMiOq9Gmn
ol7qd8bxOcO9TVXctsXgbhMsDyiOp6FvPKlCYHHjCwBSY1EQLza2liBope5ocqtAUBecxq2iUxz7
W42dzE8f1FWKnblu8iMQT1JgZtpXvoP7IQ27QYNAwLFZifADSziIQQXNDd3MLONffMCoYoiwK0UI
LeZOXBgbVGDzDDS6ss09xu2JFYqPQ7qyIXmfPQb+gpU87GbypCWGTArFZyDLoDVz9bv37MpLTeeF
jZVTS1apLvjJv+YCDAjnbiUwoKsGSUYmu7EieUUh8lGPlQJDVl/R5ax6IXZb6DdieJQpYi49xcEl
TLU3iknJZFp8fI44MXaemP6O0ydCzvnMluO97/8gd2D41rE7koukPj6W5UOHqebWHTwNO+Uxn1IP
55PSyYk3cl3c0IBxmSOx5tj0XDdkBJEtjIPLsxt7IpzctJlgvWHd0qfhJs28Agb/Sk7iTHeINRJ7
eJR6EvWVHw2xNhYp9k791WYq84q/5hoqVdAjPz+F7T+VbFdc1XLetY6yEfEsUTx/vamaw4pyDstL
4a3oirlyMOMTObnujuONJpZgCD+Ms2xF8WJ/RvyN1ijBpJTrEFnNbb/8pv3RtMBZfPelgmyRtz7k
YumYaPTOk3gS2iSwMc8ct2BKT6o4RVlKYagjmV+rH4jMWMWX5/2sv+hGu6ojxCMB/M6NUY/KQ6Mq
7k3GA45hZGCfa3cBMYjGo+EjNy7hMuBIanKmFlcPLxJ04noe0Gy3dlE03ZzyyNN40RGAnqX15+RF
GYOWP+wSCx0pv2ODK1FBgH2ICGk3WdBw6vIErSzk6HSPz0rk1hLke7IYa7ZTLZ1y06HIlmoDPQ7y
zl4RoiowB6nT0LOJHPjawGk8qrWUpkRl064sCAY=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library synplify;
use synplify.components.all;
library gw1ns;
use gw1ns.components.all;

entity Gowin_EMPU_Top is
port(
  sys_clk :  in std_logic;
  gpio :  inout std_logic_vector(15 downto 0);
  reset_n :  in std_logic);
end Gowin_EMPU_Top;
architecture beh of Gowin_EMPU_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~Gowin_EMPU.Gowin_EMPU_Top\
port(
  reset_n: in std_logic;
  sys_clk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  gpio : inout std_logic_vector(15 downto 0));
end component;
begin
GND_s5: GND
port map (
  G => GND_0);
VCC_s6: VCC
port map (
  V => VCC_0);
Gowin_EMPU_inst: \~Gowin_EMPU.Gowin_EMPU_Top\
port map(
  reset_n => reset_n,
  sys_clk => sys_clk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  gpio(15 downto 0) => gpio(15 downto 0));
end beh;
