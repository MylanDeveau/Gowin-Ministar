--
--Written by GowinSynthesis
--Product Version "GowinSynthesis V1.9.8.05"
--Tue Jul 26 15:12:09 2022

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.8.05/IDE/ipcore/gowin_empu_gw1ns4/data/gowin_empu.v"
--file1 "\C:/Gowin/Gowin_V1.9.8.05/IDE/ipcore/gowin_empu_gw1ns4/data/gowin_empu_top.v"
`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
HKnaJiPSPCDZ8phcnvrFx2l4Ui70XqfPhTaAb+wEZqnd57i7VjDfwkDhip0Ew6zIZpbaF3Lw63P5
kdOIXlc+66aAYswGkzpw5XjsEnCiDo2t1GY+ASv9Wd4oQJ8GbmPK2BaB4K9v0rjQMMca3DwnwBau
vZjyzRZ4YkUWqjCKTtRH8VsLGMiQjfN2VSa/JsWH0OiUKEg/s7sbiF/9FYbQJG3G19wZH8TWrq+o
bBHaAmQ2ZeamD/2uzCNmsSfwfaXFWrxyM4is55HH5SzKNehLyStk8PNn+im4sz/wJhWgfxrLuiJB
JFkzgee50zQk+PP0IsrMEQWM9PGwG3CP8Ml0cQ==

`protect encoding=(enctype="base64", line_length=76, bytes=162320)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
lDJbRA8OHjbCkvXIDPVNfgB3+12IvBy6w6wzeygG+JTCQROBsjtYlvzgQrbwLVpT7QJm0Rz71fay
6wWXhLSH5JXBEErjjorjlKlW6je2jiXjYppwhibn6uJ+/nOl1wlXrkN7gAyu94qpFQrC4aQTKJ5+
q4ixdt9P8819YI1kChW9VqbannqDpgDLRg4TdXyfqKumIzbFN3ca7BQFvTw9cM7HBzUWCmQPKeyR
+IbRDXGS6poFJeAajNt3IufeXJgPAsJBikEu1lzlNB8T9gkNSNOlPbBIMaNY77Iv7HEIRILGHUTI
i2nwGdx16SB239DEn06t/8IvmhfPZDSRzfZIIC98n8y8NKJzoZAT4AmDx0XBkydxD1igRIj7oimF
1jreWrOmTNPdkPa/jHd9xyZrS5vtu29XISw9mtfiIOgSRbMY/5Duiv9U9kp+KoXlUc/PNA1W8ipX
ScZz2SYo+Xi+ZsRhJ+L4s6J7X9F4Jr1+aRO/15y50VOVIKHIfMSZhc/gLnF4mdOUQ5FgtcDb/Em/
oaJMxI0XHehxCLEQsQmv8T31NaWLzWX7jTl79/eoKhb6HHOD2R4r23pbL2dlFESPb0IX9upkoj+V
pN20JXsNphiDarkSnm7XKym/FHuCF3YwqAcSwTKxecw4aGeuxvdpbamKpDTiGc4sq9e7J+05nleF
jlup+Xv/vvMA6Vmx/cZs/WHxwj9PFyaF0PkHBRAevEjB5zQXRBTS7OhdBarmuEfbo/i27+tug+Ja
QIFu8EjCCEi3YaC7bExtJ+ztSXyhAA6q4efp842n3Ce0VBtrrBiHkJQZiGqaiRCetAvxzaQ2573A
LuHhjYTFLSExdoX0wjz0pwc7bLSKRmV6LOKLarVx+9UaykBnHOVXOwjZPtyzxCms1KtbLh/EqlKI
i3lzFqf0U3+uQbrlgThWG1FIY4+cbGfwyE024iHMa2uNRUI0akDCpPG0/b7tUCz4LOD8kd2oPC08
VRrDTVp6hr8OiCwOFzWVXu5R2W8RBuAcFLsulfD+mmLrNuOSCsZpOyTnBrfIy19TLW5XD0TxbauM
pCY6K2Vb3TEqD1kvkWCVqKxLC/PMMbgJhgJ7h5x2qvGEY2cHosR71zmEG33JWTDDy/WBNZhj/Ddb
T3xZtaMQX4ErFDJjj5jLeBLLHyiU5HJ4Il6Z4FAGdowLOhkK5E+FJNzgHwvcGAtmfHUpABN8FtJW
vzldJEYXiG8PWkjAOIQbprRjU7QN2sAohWWb9kMt8UOyEbhY5Df4vTXC9pqv+V/bXpbcbsKMYtSc
UWlnEL7ZS0P37VidI7Zw/T++4TV1yCzIjdMzgvygR0myExuVFw0hpCXEVgO3R8Ub04HK0s1uZn0g
3y1k0umvaLnvAlxyZJBFe2rZcl7ZXQqdTa6UZxU4TLJzxaEcHnZ06beg5MnMzQsSEJGMiUcLxbvQ
z0KkQrxUEOfQMSNw6vrrOrxG5jhu6mObTsm8XWNOjm2CAxt9QEE1l+Wp5ZO4hu1RY6xvc5WQ4DL9
2/CXOhA1mQlK6qC+3L5GhztElUeT5c5aCPmnXmweMZND8UG7qLwllcPVshg10PzR3AjGFc6yuMpZ
1M+XPHwLKLTBE0F1MOngx+saxNL40TVnnHEz+yuaC98gHsH8MPul3YgMeUxhF1KOnbds75m/Metf
jbEDlM/AA/txBnENSUGXCx87v88EemDrZnlp5ynbJnxCegpbhKZJWEsSBUiU1AoLiEKPK7Jp0E1c
LOYVCqR+lAGILkVID8pGWc0Jv1e80xxxxxQN3UCqYwGZ6rR3jkl0hiy8QDalQ2gWmEQwOvsmXE8M
i/nwsz6QicYtxZUn4i/kFw2dFx1uIeq/wTMASbEP3R4Rv6jb/nXmL/xQH6q4h05Fvk7PglUa24C5
tW+xZyD2oGIa+4TlLi9k5PqVLvH9odcDavaXa3jmAht8u+HtP7rykFgN6NmsV8YT8XvS8yobkWZM
VsOLYoyuL5Hmc2+sFyM+YqMrhqpokxetrQd+m2Esua7T6pLh6/twNbqTdD5NVi89ZJBa1ejsRVE8
0lBA1ImufaWm+zHixh34ksyCtlhnwj+YheCwehcvcgjFYzPUU6GBSA9F87RLjXbHScwiZbyYnWqL
krIYZrPvCnbKr91VSDqM2exQ21LM3kaO10GAc7mEK+d8ofrgeqtBeclTWOHDclgi8NH0UVzaYETO
s8bG3IIV65rI+SYUCsrs+Hti2aV30ndaxneoe+xZ4B2Goy2t2xkgOUhPoSZlmzlyE3D3v+pr7XIG
/O0UdNxh5s6DiDsjMOBPgPKlfmDkMW5MM1c5rw4YiXVRzBZtdeWUKoyDK1IW2sl49ZKg4m8B9dtp
CrHDqeWwa/5HyGX+9WJeTsK60Hw6rlhQbvG2ihKGdAMgG+4LeuQm+FEmSkpmz71lNfQ8L3cmqH2M
/NOFRVZEaUzHxCcKC7wccuKJE54v02OnzS4zuFTyETWWKlNuuZiDZwbW5+zk0Q4KbhqqIXYlq2Z/
gej7CH3pgB3qTLTfl+IX4FxKBY0mBhkCiqKlwft9f7BqC9/8jCzs3FGecFmws37FhWxvxaPTyY3G
N9RuQICjpKlUs/Qi+b3DQreKHjPUIexiw2nchND9NMaLruJJ44q/KD/YA+Icvx5rWVtaGvII6t5/
OfyzEJR0gGb/5nA7iLfoxVdFXNc9kwzdD0MwPB9JJyVd/+2t1mLvRAFurkITjYvzZo+pkGJKNQfV
Zt6eVxA7mY34IBZhz0FL3lGjHG5KmogCAFofQOLOyhT0H8f7QNk3q6M8qZY6M5Y4CqpuV8ekFsgG
7KS8RfTgIWhqaKBO3T+kf0JfclhfxCKpDM/+SC60+Dzzz+hQnyA3f3Gsv3DwzWtFKyGoUITNvy4G
mOND63pds8P0xZMBpw0OsUgJNR/tJiYWkulmwcyW98YLTOG1XZTvy7GghxP6eJOASUTKizOiZSFI
2u6Ee0Of0spHEbDDg5wBkk9RDM1kLrXHc7O9Oped+osX5Yxc3+AxcULU/lOkgiqI3BVHXzXdR7E+
VkEnecHbEKG4mj7+kT+j2OOAOpNQsoa9zBzyhvHA06X3/HzsNAt9Fqyhj85AL8Mv9CLlafsOYZJF
gtDZAX1zc3Ylf92r840zG50Hjzs5MWxbJ4MX96fSAW/IUyUjnbp0jriVn+Ic04SjwJVJozC491Ld
U0dlejoleS8ujC47azGoSuV24+lh3vHkdZtjyw1nRj1DQxIKsvgttNLw8G2/ltiCoS0rCHSAZNYs
N6OC7YmgpCrqdxEYX6nBjSZFaHgG4ckFIukRnTTi6/pAjaUjXDmIrN1x8kWGzCq90m+R+inqtBnm
PwYayH90Q5oh5OoIHmcNEaKXxzZOojCdf1FMVc+iE2GFoQa+rzZz2PWRecnQFIPqmAYUl3S1z33M
0c1ybVzd30XhQ2Al5+cB2KWEb2I7rulhUaftc8gij3oebWIie/wvLIHzDyal5ubhveNCAjd1E2di
rNa58yqDrQ2I8NhnKGcChT5PIbnxg0ZQO3O2x8xt5j2bm8qKR6EzMCrQu5s08tl+0Thpnd7AdrE3
S/Sn3z8aqjOikfjiwwHn1ajcsgNhHejzoPpq59jkxjpl96qv/DXYJRbzgL3nd4hfl2uNF+DnyNyf
mq+7YPhsYgFmmKbtFlHfaGAh1te1IYRlcoABfy5qRWeQ6dOWojO0XK32OfaaJsanM4IYf01DIK2G
nhg6zJOLZnj8vsM1jAP4xkctFzjfkMieiFbMywuBLxd68rxnH2IQ/V7dLxWz/lXieIH0XhduiUEf
wdCRuNN8yAXjjQqJ+12N+HtMpw/p+7mUncDpNveTjVb/2WvqnnDYq4gbBsfGEe/0T7wT93TPVIQj
ynbbY04n4M1sqbQCoaSRQfsdTl9NKmOdOHRaxppVuMv4Y2judmaP3PHWFVzqZSG8q2xvnOOntTPV
2obaZT+T+YQVALtZJEiG80YasppKOFlhjPmUmhFn5kmGPCNBSAX5euc5Gelj0bhsC5r8zJUfM/Tp
o7la81gDXjK0plosjGXlEn0HSQEAZkviHFFIAurW+I0ObABUqZQcVYY7x/y1p4LkqTMl5X9T3lYa
7b6SBSEY76bpvAqf9SJWW9dMFiZ5i0foKgbdzHPgybUa1bTzEkuoBfqevfPWAKQ1xNkLmM7hUSoZ
Lm+dUk8/HOww/N9osUWgWuYCkwyd7lKJ3VXDZbC02AJIHGEIXgpjKvPRvK7Fz+wZZZ2BW2Phx9py
LWKFepXaCwb6/q3rs/7VmBybOnkvKWrL3AjERnOULBZFFKORaBpZy6Z00D72WKMiNvO4JJWmkGlG
8hNjI6Zu+7hnbiq6iHnU8cLdHtYZvl40tVNqzQcdIqN+IxCjUxVBEmfJPog65Wo4qrpUne2AY5MF
5GmCV5vZDs65+xuHEr7sEgaWJLUD28x1/uA0+uaFcLcngF10cdNPMYFJ4CggE9nkR6tF+Z6wXjvM
/xcLSExKqZV34U/SULXXjZmA/xe59muW+NABYdabdaVTMlQJJNI7qagQoJf77bKhIXLfTJUVdsLI
wp2r0cD4ZS/7HmY9a2yAz6zlP2G8r/9AHS9zQP19sS3A2tA9OQeCsbs5KN6E3D0sTE1ARqEcSM3J
G7ze/6qlsQdLYpzzNjh3kU2+MRHKSu9e8QIaQkvAMYGF+d/N/UtLB13VpSzbNh21sXgzTyderP3n
8P+13669yBczvXL+GRCtnmHi/q3aMcQVr/cTORi81GViPDhLfQQnxuQ4VxvXaz6j1JPBcmsojS2A
BE26R3N2RrzEYGnK9F76HoHiZIFDL/zQlCL8nCixH+4JuCvugcPrBcn1f8vrU0q6rg3wBcnHP+6C
2ipj3TSMWBL0so+AWnZeLMb5x++sPBdFkJZBL4Tbi+J7EGnNWl5gUTD1aRzpc0sAsAloVE2qFJG0
Ek/MdkqAS4mMiW4UCdCOZdZxAsGMmZdkO0NU6zlmPnxr6n2yUrFg8m6Ypu4NnJrTyycVht37FTuH
egwANZG++LLRjlZGraJJIXrqITA4CfNZf0uIcENiQwMj/sxssj8ShQNfCia/KjZ/KNDVtL+1wcTc
tqg6XzDzYHTZY4mu++q+iTlUncchlSa/kcr+S0enI73z+Izbct+FZrgkIZM3TocQO94agIQZIHoX
GTntWOJqQEFuzcSdiyQC+hDGQWiuhVq9PqPNbeDKeNUYazFDY6iJLyRM1RDFDgZSPAtqywZ3QCQy
cgj5sTyIqha7ajPZb5rsA5sH9ZfN3zTAaBKrzI1/jLvVqAZ6OmzIXN6ACiWxTu+3T5fNpzJhaudE
QB/mphGBSDTlvdhpa33XqdWrH0doW/oS0LUJhlYO1Tr+hSig/MOykvkp4bh2ke5KYauTx7/MWUTo
WcY50fXSXBG95YrsgaMDaLTw0E16bthRnYsvksyT+XNggVZopo/M1WRbQPMYZPZ5RUDxsEerXe1z
x4MSycGNcSRBplCTo2nSviyKF4c+079qyge2RJ//equSXBDmteoP+doHlkab7PesV2UHfT7BkOuD
hgK9r9uVuJXOek+KMk6UJSMOqhdO9KM5l6zVhzofOXXxSQtBVtt9ESDR0Bhn+hOfFZCFv/U7ycQR
z9DinTyTOspDm3F8plZc0eHFyoHPUZ+WRoTf22MoXQ42kwyXq4n29X0LYVXBg8GncPQ3NEOV+jiS
8MtnuSamqVZs8vqjYdGxmr6TAnKvurOsIf1lnpWMynJzbkvYYxxwAuM75h8lTB4AsKRSbIU4+x35
wOTCkMhtXo4YX6S/4LPBRW952D0Vq+V5xr+LvjktSrk1EZZaO92b2hNWDg6v+W7Ra7bRhFUQXm4k
koVb6siL9QVzfcr5YzH3e1l4kRTvh8CrGZsEJQyFfjf9XIdFK0QXKzc9AM+6ERzyuwuXdb/7IBIO
1k/ahFv5xqF2ANJSsobDAQWHHEmaoQM4+lB51NFAolXTdG9memeU9zFP01nWFcVGX6NylPnowEs2
98Q4GYjbCEGjhmw+s43Q2+g/wFWv9I9n7lgxTZG9ODm8F8Fs138KSboSK2pz2+Ki0UjbgYhHullw
+ao0jnksAB3ds3MrQ6g3ewUb6crJNISmzcxFu3Wdhf0fi6ycv6Jqd3mEf3Dh6HZfDkwOd//3Tqdo
qswcbDZBCSweSJDi+hyGgceFvW9yVshzzBAElA20Kp3KCEU+IcolDpFtgzHpHvWiHAcoxHNPIWJT
Bsdq83IGtxC16e8IIexDGOD3BdMf+imx4njfjMiStm6GbWDvRzvSn7S4cPSKlTRMkKPvY0lcamEf
fR2w9w111FZu+zdakGn0KnUkWXfBoyEM2bEVwBIBYgdtY0COlcavfg+zahoZzykiMyWio7OnGAo6
pccCNlSbPziXtbhv/QCLywpYV+J7pO8ZArCxg9qgBde92nvGSFlU+JhqzvkTxHCZ5JMhpA7kZO1l
cam5yelB4mU/AEMCZL5Nk3FXTJR1CbaJzdQy4+wBynp1Hq+tVWLFi8gHTTOTEdVRdmXK3YAq0Pb/
MOj1H+2kchTxU2dSmaA/YBckAN3AXGHd6eYjp7AtBekGI09k7vOgNBbVily1cA18aMhDdJuZ63tK
bemfmBt+VkLzTEdD8DkSiTkSFQJRPVnDj1r3bAEGrsyOtTjtG1Neo+hzUygqjD3fuB2A2Gp+yHdj
mJrsi0kT+Rr5BbFKlZhg3MT+jr6l2KYyEiM6IvpFCqhVY8jcaQ4w1tFjYxgJaEeIWERIGdDQGsAk
AOr4qojYmi2KmadiOUfNx7bpPAszUJOJQEkY90GRLXmx3GuFSS8CanhX4CxCX596wVD/jSRxvsSQ
PZB9sG5GkLHOYZezPuiMFYvpsQrzkzoOLBg6sWrcdUqbWN2/qT5Q4FIWDmqYLNtozuhbBk6rorku
VkYgV3rAcpTVGeaUXImZrCzlGNgQsYj4mrTKNmgr+5LQzJm72c1rPQDcAKhNScbyxzinM3NWHXg6
ZsxQY9kQIRQ2TIMkyVSHRevxxT5TxIq68gFzhJ7+QF/weDzDln5cMXmVBe5OPDhNTb0fMNLJAXUM
1tUW6caOflDH8ugOrWGd6+nF8qG+KclbH3Fz71G5JhV+Wp5GdPvcGQP+gH3nEni9V18MqIeOcKRR
PT4gw/FYlz8D1R/H0T9n5pbgmq9qr3DA5ud/uZXZ/RHnz9hSoeqi++NNtFTAbrFdDiqD2VEZkV66
F1xZ2vxgC3Fdd9u8ckv2zMyWPGfAko2PLWNON0YM/p1DqhFwjv4VJQkxgLKcqXQNO2UXAsJkdri0
zGVDO4TAJVBmriyVpVwaupoG7IFYPy/44JW+sLzMqfRBqfjgeKsGidNhDxYf/89pFLBLQbzi3pUE
Bs85+mSBrPQWT1ymxQe/dWWK2OD2/GJX33/O+T2Y1SVGzWy3VUG11Z9QkqBiqe1qlRUdMRbCRI8O
aM3fyPu17X1n8XzHa5ziIfIFws03VhcqOTu5DJXvTvu7ta5f3UMA+ScGpRM4THQXFEkbkJVFEceI
LRZn+pyOhtsPA4FCdjZnL/AXncG1hdd8fOnjPNOoj2wdHmDOsa2BKpqChWEnNjX1a30+oSKHPGU8
W+J56IVemtrZB1//vPN/7cJNOSc0B6gCVbeG9QHV9BWsB3KynU959Ruas1U5SvZUZMBZMInUjQcI
fwTIhbbIS7rIFHcf+P7ARyG8ciUYnGN+0NZgvIvzfASFo8wJrb6JMn1brlARakuvn3C2/03a5rZK
J0ACfEed3ge58uxC+dN7qcnJaGaHeqhhpZnhgSMq7yv2ZErhdQY8mfzVzzE3c2KS3VdvQfugqegx
urWJ1g7ZqHIEjykVvnRE9pHoKo0S/dHHJKQSWHCLzA5W+VdmgGLcDBGjUK2aSz1ikrIHrUfVBx9h
FqAr9MEDhPX82R0KL8SRpXe7NoYQCg8gOqgj8nM7eqfRRM0vJ+vSZqhVnJbhrkbDTAwo5JrrMx8X
PaJxaUKtp7BSwj8S4NEN1fYDDjyCoeqU4b/iVD1jrtAH1IclemfFHBFam3OW2eFEGqjXowtHcfpA
5thPYSdqNM2G/14n4GHHo013HtW2uEy2rgTt+4dy48db8EoRxafXEnKJzsy2/poe8zHBktv+cG/a
v7k6B0V3yeogdUAHo76L/N++IJG0ijfwiVjW5iOL7QnMTcBvkI1vYdTor/zGw4Xc+PG5hk1ctKnk
39uw1JDGv14GVjfqOsTrhIyAP+sPM7HsieO7RyCadvxqZik++Zpg2gwgmt+Zzp9vgM4xsyayVcMR
LjgKEw1lg/U6O+dW3aFfYRldPuBZu+/TvTbjIdTDr26xp3jiD50CdXnoN7q99akvSi9vKNTkllhA
z/dCqAGGMNXgguOIjti19Ip21fRrPnkyzuNVC1ezTT6UGm21KOx1W2fHMNhrqf7wPhnJeY8dRHqM
odl8T+VH4cEvFGREPH73xUJvWjs3hQWbqKnfo42Qw5m4mffH75nl5FIKhb/wtCYe/hVhW6CUcfWw
/OzQktgep2YDZzriGXz8UfB74mCNE0Ni0ddKQoO/EteM4RW23m2G553LyVvyAqHULm7AVFx/db7d
XL9wLN1s23vj6yA9cmPQLFstD9EnU2plO2z2V1UvfCH6Q6lpjz9PQYNu/1aSWOmwUger63fNxrGl
rxIjIQW6pQsF8g90vE6yJvffE9gvRDQhYbt4o/5sT53s0Ni1nBhOtTH7hGOFaBOfchhwceIWfEIF
WLU9Q1m8XXZxyAkM3Aj5XY4b4ViZoc5ZjQF1iVMGvo1OWjpPxrbv47/AhrPNILiQWO8eVilN2hw3
iW2vH1XwI+aDqjdBDNi953sATu7dGlk4ySL+3q5GyIvPWhYO/p37Fqum6fuNKaCTAa8iL/sNb50y
cySGqQYpDvZ1CnJ6Owi9van6WqLSrneydQPmYSqu3AhHKIcG2g7Taq6CBVpvAsPROLmRhW5BzYVx
262A+R72/N5r8ySzCwqZ92fwOEU9ZwvUkCk5RJk/br9usAMJz/lZ/VyFsSJ4yMRgNfXFxgJ10MHg
XnJF1n4fz+LMTpAcU6C705Mde0gcxPMgGLGDSUizk0UtmhP2nBRx2HW2a9Gxu6IyNY8+JUfkW3ON
ct2Ef1tiJLKzG7INP6zxpwvtcIi4r5fAOrA8vNbaWvX/JB400EvKvjH4em1VroYIo36Zr4PscFOr
3+zuxQ5sIqFBbty6UCZrjWKJZWNN1a7J1OPLFZdi/WuJjZ3bGKWHcmoSSQrtSD8pEivXqhrWfpx/
tcKb58mTnc9v3Wpta/QZLqMMOod4J0YULy1mxY9CZyBDmqspjpyJogdUFC9ITA1E4cFoEKI6tDxk
009CGiB4ijV/l8RNsmJvdPrKhfN+DTXmSOro/iPtaoAuQf1bsPJ6+mEZCQAwLbxZwD4O8Z5+FOhZ
CoPO6N216EF+kGK71PUp0PGiGj1abpOMasEeNvdgnTObWEwg9l3SZh40xMEHsUzI5/q0FzU7/PlD
YLbXwDvfEw0hamy+BDicf6q0zsk7tu2vTi7+fiGnaXaod9JlaiSSoK85CRE0Ev83JAQ7LeiRp2ob
cDFnbjK6CFWftr7MRJ3jNu3hEnudYch/pdUAg46r+S+oIYQWBl4U0dCGft+z7stabWO7Q2cautBQ
IgrMyoTjI7rVooBEEuunGcj13q/wVgFd+YfRf0Sw+sg+ZgHTDF3RJFZ83DOAtQ5ncr/KYz18B7/9
9h1kaiQB+4t9imUxGDHlyaVJQeXs5deFfEdmfYGsbyb/Aza7+Fn8ZVhLHNDzIe3BO8t+sXHGepGY
vwhHMCzTui6T8J3NOPFbD2Ejm6b4s/tvYXI+NkICDwL/wD762MiZat9Q97oYap1zdZoPEt7CLmR4
8iDSzwv4wjQlhyiHQDYssGPW7LXgXZAZcrm6negnlzv2dXap7eCv3Q3k4Wh3KiMerJXLgSle7T9a
7CHyCTM5Dq8hDPkbHxuDhTXy2S1xaIeEbUvm5EUJqpzoV9fhn6LvPZe3jtAsNFU3YWQfvHO/wPXy
u13eNropukaNnR4ySc+A3VD8RhyHkf/4AohIJgMBSqTg3wF7XBeV7Ofuv1IzptizyHL3mpwQr0GV
U2YWbvePXDhKtqNGeEPpnix8L0pP7aSQeO4/hntOh4BXCXPIxc4l7BzlsGYOGGcqk2dzWQcFvWv9
lqsVKeo9osnAcrnBLPWW0Smj022edfqiysTq1VQELBgS8R5CaTTjuhgSS16mvT1Tmyzas+6L47Dv
55SdQYo18Z0QoR7P0Em/ixnKRto7AYU+XIjCDFJRITC0x6ZDMpRZNJjB3/yr8wfD3A6Td42bh8A7
wFuuGXnAoAsmkjaPuNF/q0Mpb8kpaNbYIhR/8WEK3PYlX4kBb+PV5nDru1b1i2+6ReGFGdnZcZsg
PC9784TUAE4W7DKUNtxJezXF/NNQGfQ6/Os2fmUqqTQFykv5mRdZ7fjw1VM8P9jcFSx8wjz5yyZ7
DN7bDuvsVjmsqRIPNEIqC9Zk7wy7EHOpTP5KRLxKfz5t89rTLKCfEYf/tb9trBaZ9+YVFYasjd1p
nGcY2qM4CyK4J+tmIsqkn2wZe4vAfS4khc4f+IHSLzrMDrgtc1heC21dR2MICpG/Qb7pd+OmO6uJ
PFu/cRo1EnqnEW7XLnigBvBxX0bW3CRGEO9VlC4BuHrtY9aU/g/OsdlNm7TNVBhZpt0u5ijZ4vV1
8oHsz3brH3/3nI/9YFEax4Y9belTE93j0dtW7x9OTTHeXAhRwvLc09AAemTV1jKsWy8T6fyJHi7S
o58lFSHQnm2VtVSjFIjDA17qfafGAQmpElyzhLXUaAVJepbwKjhFJ2NtG6nJz7E+Z5C3QxVMyJdJ
+hsNNwnS0mdqCrCA3u8pYZFWpz7BfamPOE7eLEcqZOMAogZUNhXSvBEvX6fnBVYmSUtNLvJu7WLA
r1KpzFF2idAomIKdbho8HNGD1b5Em4HnrvoDLpBstDPbglXtJ6I5mvYJiWB0x7IZj+D6zyT1Felr
yp9e4jZrJ4Mxarttm7GH8a8V47xgJfJ9B/v6dv2SVgHPq++ywhKAsdqVdNyHPi4hlHRCMbvMRo4o
UXqcSNKbYAUd5PW78gPhzxwvxKh/ZJMl/7NkubHqgfo5uUbLHn7LRiVrAKasXpA9XuPq4M3Q0grS
kY7hlx1W3p8kbyrDMF0EA58ujBOsN/XlsTKvl6oLPaUjTE24sMx1tITPHlvHapb/qin338Qa7fzt
64tHXkhCNQ1xEKOQ2qqyhDMYTQGMAWZydJmUZwxhPpBxOM1s4Zlz7VjaZgZW21sByHss9RlaN9H0
kvz7WSWhJiQs55DRkb/J6IOhypR3RWzcQ8qenK/6WqDrXfMG/d+5au0qtUt8dQqp+aLw5oF20hxC
LXM0z4zZLQdY5XncA3R9qO0GlaSyxVPq3dA4KsptgnS88m0eRAQ2yPokVYHAogcLtFkUrg/2O+hJ
6ks0hIfLtAEGay4vxWjp35IOFZJPpgyI4VHnImgOO+1lw2y4VE33AZGaSFw3Mt8YX6x+SY7iEP5I
i9PiZ/lCUtq+eTxHqX+UO6In+tYP3mt+9msISzccRZ/fbiCGkx0rmdsKr3+ZUaG9+xnvz5hZtpuT
ZbUv0Cv2it+Z5BJZ3khpbpZqgId5mdspQE4rkLRr/v5wedp4N6ikEMQefPC7TXgsSjr89UrvtRKU
135cw+uO+QmYYVkJqNUgMx25Ene48A+VV4uKoz5tOMvjRUg64b9kDfm/1PZxtdriKzsHAMtuaeSJ
BT8XqSsok1Ofsxv3T1rfCtPfRetI5+vXvV1Z4FQFM5xpI2WVuvEBGftp+JUs9lpX7d3UrO4Vcljr
eZZmipRa7q7BM61sXoAMZxBmKDfAM43pzoZZ/hCgcIfVMeMG2vOpVWubsNIQVz47XvCV3RBF9WcA
mVU9ILfonwtM5DgpgW+1p5MxuLicN+Fv7scY/QLCeu0ZYXc/Z/nBvmJomOuhFLRciE28EE0vyurl
flcMkg+nGUXUrv0HyuP+0+tZK9o04Dn/JTEcDavBwBPIsNx0FC9S8p7FOOAtHHdhXJL3DTZFo19l
0Bbdi27ERJNpVWjHuI8GWQ73cgAIjedyUvwg07CJCeALxXiWi7StW7vYqwvGRIgcLbWk7xJsL4s3
M99gzE6VZZHdCOqRIbSv9RMtyoIKR/IaRRAobINYOtd4R5qRkaR0jrQoBiAo3w94gx52FTN3Hi27
CtuoAzI2SKRCHmRFfWWaf94+qVHqLuwMZiJTVRqSwP5ZWLbzoHeib2jK+u/1huQ81C5125yjTZpb
b/71cu3cZZvum87iF4SR41yCD4fqgCfNgiw+DBRWzTjVQRSXvs6O7tpcf851jweaEPZhoj3739JP
+fGnigZPkW8cI/rtKVW6ZrKmPRPxDC9SuCuxrEnqgWB1ensV1OdLznQi7Db09urOmY4BkItWbRX4
NpCy12IznANdVD2TsT6v280Pi1Pu0CoxmvwbK461NGwYsAmRkXusrbIAXv0G1eT6PfIIwJrbBx6y
icyLcigLfIEL7aGFeZJyCPTuEAhtQwQ4jMXgvg4gksDjh4Py3mBHFKK32euoA/Ir7M4OOnGCKQ1I
H6UGZF0mmlVEyeyMgUIv0ciORbopNJa32w+FZMUdcuB8k/Y8gKVOAKc0pYXPjHZGJE7phc/3KaUA
97e/mNoIM01W+1cwds70F6PufJcpbHMCIjNsGkAB3n2YWLBecVzheCwNe3fiY0fPO4DBG/tGmY9y
QCY6ew0AJBqhr4Xkn8wmZFRUAnWNPa0u7HP8oH9g6zcXTBDlnj6bCudefOxmHFEwn/7dT2+ny/cU
Y2hnICJJvK6DUELbBe1fQBtghRP6Ft66vFVLEB/jb6xEmY1fyKAdtswppv47qvWtMxiXlU20ttKn
arMiWpGGArkT9PjPw9EAGsrlNzMdWGrkF5McoHGHcXwKTZyzWsp67TV1ho987kuxZTphZ1o4G7vs
FY1y6u57s1nAxK8QUPm+8961P5cX1sOPVcmyykGAhDbyobCfE75PZ9yDvknjeKnHDoXg5xXVlcxF
mZWOROU6licqxBVjlR3Pask8sr/V5m6JhVcmH6HE3sa02dob5Rp3Klw6b9Op3xWm6BNcijd/AyNg
0ZUDKb/azXyq+saHVBiyQhc4ULbH+Fv9nQPc7woC0+PacUYHacOxkdwXWrVH+TO1td44Ran0xK1j
t16R7NqYZzg6/tAc5kRmdph5R//f2nHhs/tZGfL1VzyO+/PohkzwTF9+eNYPss4uc6niL0lATtkE
AXpxFgcoEkVgXXSx60vpQCzfNRk9/MnNZzv9MuXSHF+F51XHu9n7lcOb5iFWUJrPaxGLqkcnQM3T
SHKjiKlwgmZdLbuxRZhewi03hE66vPxEi5uZqJJW5YeqqK490qzYGNMCfK+pAotUqkb4NqMklzIT
HKAR/H3k5wzQUr6SJI+AXCttWjzUJ2dahjVR5My76cwcW5hiKSiRrFQ0n/bMTog3ctZXZBVGgvij
BGGDgE4LBmfjbWQo6J7oMEvuOG3WAYvC0AnJUfmOVsWqBz8CVeBiE7obz60BK+CoH3nS3BvfTDWO
wDyWV2KFGPo9QyZaEjr9CRqdDt9QEj/KnNsOW9g7Gi67RpiGs3O7iKOhc3tTSuHiC7A3xjIkThua
4hBOoOSqwQgTJvOtJ8arM4KK9c2EDkIHEaAxHqAnVKHs29pe1CXIz6k40NCZhFRpE1nHY+fjGsaH
4KEvlgBrCe0yTutgefCzPxorSpFk18kUEi0Ca0Wh3KRVZKG7Ty89cc1Nr1VvA7ubsVTzWx4emU7k
5N3fKzkbQY4Rt3O0t3ulzJlP57FoijHPA9K/ScfocWz+AOaeqM9AudGdXeheMqLhpqsPFNQjhw1Z
IYxmeSG2R9kHs8CI116ZqcVBlvy9Lg9C2aD23Tb8e9UySHDo55FkSz2VULhjDOhlAgrVhy+Y3AOe
laObR5YT63Jy/tmj+f/1Wg3MbhYtfKSKQXj56V9lFR2w1jtc5RPDWd2Yein//OOYODX9BlIn7gJP
lZFp6RC1kFeyZdhx577Av9EtUMy9Djb0RGsdMIS/TN10Vs5GlnfrDO1gdm6EZzbKSRjRWK1kdEVw
NgnmOLNfQNwchhAVKj6ZuttgOF1PZ04BfTQQ5G3Vub4iS+bqRW8Vk9natw7F6FUXw14/iyNBD9qW
Fu1CxlytS/Br4ftBeJ9qiwcH/NEL5dkgI6jjxf53lASvRE7Wo15Nzy1kAilOWd2BCVEoJKap6e7g
8v2jUzBNS2iZL7VUEr835f9EYnx6SqUzdWDnrThZyjFTkdjSb5kT3V8S8mLLKJQV3sSAFLghHc5z
GCt/yuWVUJZ6/71YdWvzTKf74wBdoWF1EcBlqX+MQs2sO0CwVboydcLM3ot1zielF4rPF8uJQE8D
JQQZT30tnTHuHptjrpBjgMWioSnLpXK0PjyS723qaHTOgqbqUfM07624KpDPBZLw99Wqa5r9JnBN
FIduk327lMJmF2CxyHY77QTtQsKZJHqIv0r+huQGAjzXvEkD4VpvUBLVv4TWENXIvBsPcXLcXgVz
povUd2YwCRQt4G7orWAT7wGJwVw9INJgfU7mLZ9lx8ezZbPhIMR7ewDs1e94fEQOwbAJ2atcptXt
HaI/JHOwVL9WjSAvpWr1irUMW6t6XheTpzJhIOpxm29q8Yz+/qam5Y1feWS8liAPQfFXRvK7bEJw
dwN3Q3qELp82LHtLMvODy9ya4Fn9SCEVjH+Dqx6zzEk79efhv7sW+y2mWBtaWjbTEt3J8VeSgy0U
0kBOZOWMsxytSwof8khL+ZNX7apvVKjgUSikgtUaPWcdcvof843M7HwcqQggGh8Mf/q2egWYr+Z6
2VMyQ9wBQIx+DOUceMr2avFWnFPshP+asjzlhi+r6hpNVRu06qaGeL+FO3zmEBxxgXbZe2ie0Wk7
HVX3Llj7QaYxy9wLybUZUt3MJgypQ49qVYmHHcE2eja2DjgN6j0FMlrPpCYnXGtKzEbLSsbi6gBP
ReFHOlwOMhT/z705xSv3AqFQG8Amxh8hdQeZSzXxDMFzzezzGQHgtwQngodeGT0zZvNUBZjTm1xd
eaIblZYhl10FpyOVFeuCVVg2rs9YaRpJIhBKVX0L4pUu790Xdxj+N8KuJShg6WdreTlg5XuUaBZk
uAsNPBUu5i/pP6O2p60VUxPxZHHFkOqTl7ccld2bhZjjV7DFokZJAmSOYS0q8Kl4Ep4tTFSlelDR
vd1a4AMZmj6qxMHbpe2vzpQp/OMHeeLe2BgApvFBHASC9wDCsd02pzzNHQgPYUAJ4igLfWMYY0Hi
wDN8B8Lo4U1XSTa1fdQvCive8d5fqp9nb6/FjfF02mV/dJFcwuCLAiW6EnI2Yu9gAWSVkc8Q+jf9
o3ukoavhb0xoEIMRXybSCANNQqqL0vUPNl5RWWvPCScKjVdyJ+XbwjfhfxZPj2dwr5cOe1WFi8/b
HLl+EXrlCnm4ttiZZD0Zq1AFPK6evWqy2VMbzl35g8PuJ2LEQODSIRwd0xDTANf21Dv3S5G/FXiI
La7rCmSa8VMHa42zMGsjISANo9Y6oZpLRmEdVuNPnAx8r5b0wSn/928zU+J6rc6lH/pToCOtTrT5
4EZLi8ntcc63Zywn3jo4+67EwlyMxqFnHs77EQ7Ia36PQbO55usLB1OmAg1uDamNLa/dd+NmSFa0
Q0Tf29k+xJSneeHKctir2iki8mpyovEqW1BhDaTnFPnmgPaE8/6cnglBhvtrhD/qqZo2VNsusN3W
Yf+bXp2Z/f2vV7VwS7XE9yMCZ23ODFvg3nY+Dr1Yh1kU0IKPg30xg6mvYidafQSSqhVOV2Y9V0Dl
z8UbB9upD/LwUwvnT/XkOMhZYmr5te31qvPWbZIPI831iuGhpqOTYpYwMs7t/Z29CEt9r7r3BnMS
UWN9UyfRHSs599KlDOXqYf1Ypj0t8VO29aiATIIqzbAYm8muBF6UaZVVgbJqz32DX2Wf9Mn3RkZ1
MwY4+99pMoHf68SlUoqd/xAMZijRr+N7hTExmqRg1olS5AcqsvbOjiqaGtjyb82dgVqM4ddB36dn
bLfDif9XBb4JO+sA6IpNjpu0nes4K7w/GHv4qsPg0YVybOeXy2Ezmu54nHVmuy3zqsD4SvME6FGG
lOKSR3S6/pa5S96HN2vfsKXzK9RHUwOaeTEtoXIkit5MR2gxt4HRt1ZTFGBPYxogATTiYfmYVt38
fHEWYJi0ynY7DdJJBqvX/nX1RF1LM28zjGFaOGykd+FzgkV12IJVY1FwsoPUldvhNH66fkK9ATNa
wwdOQh7E91SBG0Ag6aGkgPojgrqxvpgtITe1YIiwR8UirqmANZJu6oTFj0Xel7l+a5AgG4p4ASAk
NS3C8jRgS1aUaNpQAS2Jl1OZFD2wpBd1hYgSVN9EJXjrvJp2VFFB9MBegC9hzzc1ov5OHXJ7/GRk
jD9hJr6kcvfbWQwlZMguXh43BUj4LIJb8p6kKSpfRpBM4np0bgbLsGZ/IZu16kpnWLnNQ6Wn+St/
zVvh0YIS5W0ZVwyJbvFX7J9ShPmYjj/aHKtU+N/3S/LFZZm1XlBriSxQA1lGB3brnQh5O6UFgokN
x/eC3DPsfZL9NwWtTCUz86cfjL65y+KSXtG/Q0C44RWmIjluOHR0zDnCoR71SbKkeh5SRR99o3Qs
H50TBUtDh0VDWolN8LycR2INei4otkTd8PM8N8y4T7or7Z/ZSsjPX2xlveK7PF9CjQEnm143dniC
w++a4PIyXBZH2LnTiyYw1UI3BlXFCVC5J7DrhvhvPU2bBuCsDURHHqqXUn5kWrIiSfJp5AndEzFp
iMsj1RjMLQKg2NuxRX5Kx8PQCZCbXI4NYGEkcyfgee/Xvo0YJRFrBkPjtLtyQBXKO5JizzsI6fA2
x51xiP1iFjv4cb+icqPhVHBceoZAgwDqRDyNX0Lgtb0kbLPYTnoFPojUPLJYVIDlkP1NmLg7kt7G
AfZIwTnPHgdZ7HPG1QbcT4DEoFfEVvr69OhT5pQpo8MHpXOGH9ya2BfGqNmrNhQmZa/xRfA0edYz
LdXpNxl9gp9qehRbMrm75CP6NtgerbzbkKY5H9iEetDatKfbxRPqU+ITUoPhz4yJJDZaiJGbfeSm
KKAPkUPz+ePHGHCbNzA6p86SGUcWGg+2KE+ev4ZqsoU3VNJ+jvi81ulZe2bRn3xvVBoqhb2Bmp5y
Qoty9lF9Jzcb/PaQYXjuAV+kBqp65fKvFfsa2TFb0lcHI87Kbkksbdt6/HPrhl7Lb8I3vmxhKr6K
41TlNM79QePVjCVa4GokKx2XamcF6Hb4QjbK5ERsS+nDMK//xkH1dJzv5QPo1y6FSX64VcS5O+fi
MbmDhktiFXv0l+9/ShjQUmx27xeeTIczTdpgzvYJVvzGJJreKaGOMiSPfpSuyBcTkOxwBtNnvCqa
xJT9wS7PMKqs0nWCtXQ1CtVsceVowjlSZ1vbre0NnugrWJtAsfdG/K75kEDDEGBb/vQaZVeQ8XmK
Alp/D7yvdMkAPUzkBrXBHyTe/tX4rYR1e2jdI5AwbJoUVuctMC+eqfFoWaRRRTbFwAxbOk6iLE3k
a+v4i2hNRwqf3xoJ77nlLG/EJuCIjA1OxedOpuaKdOVb5sHAJ+91FF9WJpCZjgS0C8i0Or+PpZJl
WtipsX77UD7sJC8vQ0wF131/Hd/nBbS/mQRiImU37GUQKHp3LMYTifhX2MG/9bgk2bNzquCEPIze
PUZ9ZglzIaZ3Nqq3gvs1/0zm5My36F0rakXVozcfU1vEY4GcIud9mFIZPmLE5IiVbnlaJlC862jv
ddl2J0ZuFwwjyZSsnLhOOw/E1IabeTA0QH7qgI7ZGwZah/llOigyT1hO2gL4PzaEw85I+VrF97Jy
Msx6OYXjhEXp9/P8IcvNsTcu9DaV5SF3aJ2dVHPLUyAmZ2zFzcB8bxg6K97hQbSbNckEybi6uuJr
xQ/eRWG9ruPVBniMio7HJOIR7Qv99jr7gKaa3KDq446wmBpa+suf6B01LeYE4OpCH605KtS5HrV0
CsABATzgBa6FUXHUYNH9H+1lzxDPS0jPjyQiZz7R9AAbFhECV3Fh7hEGAu8iEJtgOkEng/gOXWx+
roCfwDy+bAgQLR42kzxjAgffCNCRkcFHldcKtb9R+MIv0FKsqPVyHCNO2Rf2BHxpJX0qB+CTtQTO
J3RRlxVgo/RVpovntgMLUBX8XFWyVxEltSvcmzsA1tD++ypjJcpZmebpWyjXGlln2vAapHJbBb08
9C0X+L3rCv8qozl/qY0Z05sk2rsT6f9IDqTtgLStVunI4dVIuPPmO6/6wvvFgz4kyv3kxCyYyYky
/3HekPwJbYGaTnQpX4y8t0iF3/t+BY5OOZSGvLSBy/kAaZV/L/39Wu3ybojwZwMr/Q0uF+k09vAB
8/8lrDrzgu364x+evoNuqJsRJz6IxkB7fpIyF83F5m+Ty1ncRrLbuiC6qVSQ19mA5jFOYTMoO2UI
ukuFNQEl9qD1/s5NvWgWWsNGbdEj/1gb66IYfbzvBnFEWmv9xkDLKwYQB7onuziTlX4cR4DMQadn
qqB7hrMSfnCLlHGmfoqGAR7YoVVA4qGwd+pH39xrrVUkVnGBtaIb79td1WxlkT1k9a0+S4RqFby/
2D5BymUEl6JgjuHTXJw5/IrxLOZzWY5ig1UhYVwOhbfaxddurkLY/BmdK8Mve3aPudf0hiLnaqJL
k+r4pRr5/FIPQmGzrANMlNfVrx5EWvJ9twl+ZIEA2D2w79zpMFKiGSxr/1LXjqeVhDmhUGrftFbb
Ksi772cIYx+ns3Y3jKaNW/dvRCiMUw8Qjeo1iZ45+3DelOEaVgtbD9V6W6YznaxJMrAhOEDjMiX9
J9j4d7uaUpHPIdY+BsbUYclK/NCob2kRfAFKZ4bIjydPJvjiyLLTArx0ncdgUKS0tVZfLXlOkxId
FfTPE1/bQ/rBTUDs6Rtcpy3Q20S/ce3PIQJtxoKW8tQEahnm8HDSVi+5v/gTbgfcEKUqfnsSFDRr
4XHRtZ5FJax6jW0gFv+c4huJLRvP1Q0bsg8W4d+tqi0+lrs3HAZNHAGPixC85lR6H/IZTqQ7MUcT
yuj/+ShzQKwxMPDnoReB5ebsNXk0HRvrODZwRgkod5B4Da8eVjlh5wYyOMpfX0hQ0f49cQg5fm5d
oCUdMO10WSMl8Cyve5UYyCHcwv/fV5LN7S+wwhHLYNfL1G/HE6O2bWU4Ou6rJWp8GhvZAli8nvlf
Hcuo+6apNmrunsRDmUgg3cRQEgEpbY90nq6AY52uno+HIHsU+N5SneP0H2s61s10ItpUfiwTUeQF
XpGoeVY1Zt2xE2uVco5LwH/bjoQrFdrhUDDVJoYXayhkwuGCQ5x86ZAfT98iYei42KEx8fVsF8W9
19W2zxw/MpN/DfZ76qHhYf9yvBielcg07L/MXfi4rrLqBND+8JznvGp9MFwqUSd97uUJD3nAs35Z
B4fEzlYk4t3bGJAV80ka9nCZInpUItZygyb2buqclk9J0fhZuuyaQI6kZy2m4UZG2/zTfc/UIA16
yW5KM4YSvYmIBvQ2wCvWj2Wj+msZAyCdJ4CTYlXyO9JdCSRaKPKGsVZ3NgecqF9aA7F7xX04z6KM
nunske++cXjjIFYspfoFvggTf9i6ED8knLwwcoQwdG5BZSelj5daIRMA/T5tW9b6VhSOi7w3pNBQ
vFoigkTEvmxkuCCrFcqDimVL/zecNptLMzrKYGDjDRMMvMNFjYeiLP95BJ2lEpC3kzu/CMV5ECWG
plraB3oSBfY6JBLfAe9QDDanc1FEzn8WG/+SuHKlGob6pgSs8vVbi0nWun6HeKgSaSsN0j2t1FTX
s0k/e1xu24f42vZ/DcZ3eWyEAZBYie+1mGxCmv8xvOjM04FpdCjVpgVUeOU/6xf5uLBu6T5a76MH
JlFLaxutI2gBFpjsGrd2CHBCQ8yRggPDmE6kJKxogA8lF1DN1lxupYXYgLh3gR3calcV+tgYca3S
jDHbYasa2vVLXlRYxWQAuDpDnguSK1wjfaOP5/bx5bMtmct2X0lmVOGxoTl4zQHAwvJ09GMpPmP+
FcC70tlDN7WcaAfQTcy+WeMdGUvPzKgFemvDecD/KN45pZpRLg6jTS6b/74J4j4PKv4s+p6IHFEI
d+dmAxw3kHWnXn/nG52ByYpiVxEqv2n6Op/+rlDsbAcAJArB4c9AQuBMoMcjCjV5vr5WnlgC7hAd
LRyAu42ysLnixh4fM3nm3TofSHIY4mLt4n30zDrdvYiScpFfxHbVOFmXHN8RXQxuSenZGv3WKvVY
KUGGto5xs9da/oHhuhKGxpMoYuysyiRB1pmnD7nVYhQ8LZ6DFxI8tK3kGZCNN9KyV6u2BOYhdzQa
Qdz/G9AgF1IktgkACDtI6T5QJ70H/axTAM6NqW0jEFxXRylTUaIDEdToI+veGD4wYbATpS6kB2Ww
2ggPo1lV86OxPqncLAIOXHj9PzCVaUR0Zl1vm2/Ll0+/cIBYSrKbDEenX+DaKgwfLODNdehFaWP3
pnDxnncKwjNF0q7e9gTftf/qYNtmf3PGZ7PwnJensYpC6sJj/KeUEwiWjIbLnS3C6FcbyRxLWU4S
uouSr0o7JVHL2Qr1JFkotThMgUZMEaBBIOgZZm4uY9FVFN+g+NAWFRVD/l/YlVuIGSOL/M7MYAMk
gUzxu9sKrKQTLXKjpAWMGmh383lAj+gibJUt7olEbAGKo1Ko51eDjkQdFVv54Aq3VVAYy4fsqfg1
SqnN0aQTEOulH+AXS441kOiC+gxKT25upFFGbOo8W53W7Wa3PzJJgKppfVVcxYpJrFUjZxLL+i3r
YFnq+fxRDmxs/oz8cpQl4G5D7W8f+kWbkWWEjWrCWMSa3twyhF2n75PoHSG2bzBW+Z7DgXv61Zg4
mF/fhPqBcKktrgUvi7mxy13Yeko7XNKmHNJbEhY/5q2fIzbQZ49fY/rdxLL/ZIu/zy18H9tWY7Rj
9xIe6wfYucGe5g0nzR+zs++/HUxMcH9anZV34m5LsMlAYMlru94oUiSSCGajy0xm+YX3MtLV6qnu
rPkYBqZZIpI93eHOGAh4CrmLinWdiOnFGugOfP4+z2v0SB+7D35okUhtV1HTVfCURJNulbDIQMW6
0iPN14PP0HzpojK/yJn56r/7fig6N8tcDZgqM1eZFcbZopffECCspkSmh5CtwC2PPcUIbCYrWdBi
a5oHQc0BtE6ar13rnmD9sUAQbkQ/WBHc7lbRCJ9Sz2Gdh+2uBiefl0fXnexczzGsPGB4szlnAixK
WOpYsVnetibepXl6tvfaGq0QULGDYo9tOmpJnMvX9SGlTww/BMr0fRRrZDSvL2YweNFO+u62JJqI
w1j6RilDPBSl/RGQ3Ay87Xnjx7Bel8l8rLtEDfk7gqX7PBvH21roIXmBybPC3Et2zCloDJdXxcuO
2I9amEuj5rDx0g/rHFefnpgs0dcsvr4kz8KytXG8OH0CmIDLua3sHqEJ8K1NAMWZ64Rf83mP1YWK
Zqh74mmDbkF1YTJRj0dUKgmG2ZT+DDt6MfsAXQngcqXfqm1cDfGDJEjCJ4F+tjDfxDUeUvFKjlm4
QF7nB4mmuX2So8zKBnrd1T8DJylmUzPuz6RioT024U3iyi8iloCqQWVG0l9KeM2KAMoSjAl+9NJ0
MHmHF4AIRLk23U4Wxr5j0Pkw4YNxWPT1AbHWdEFPXTEbwbCWVcPZ7ICYf+O3tLiocA4yyTCGmc6M
oTpYMzSJu1dzr5N6RtwPQL2FaMNqZy5FBI2ES8FeswEr9iMPIvqFUDz0sxj9mo3Jk2iXXu2J7B4N
rmDYxgdEFdKwZM1BNsTJL3SckN8M2TRUTC1BVNtoxOFMgBqpdIW3E6WQcRzTrYft+FwC0wl37IUP
X2HgUKLHdCWTFtmJItYdO10fGay/HDH/Wuw9jbVq8VSgA8Sl6TlaiGm3rcG3l/O3Fne0StK3K2Bc
A0GBkH5lp9hADB3duosweglg7dB93+uICHpckNnW3LczN3afEuj7eecMFhhySNUxJ+BmXS0Bw4vr
VM4CkhxFZCxYWaDXQrCbyPxNLKOtHzXkjxJv8pD0xA7dBhSzuYV8SA6x6IBZ4q6flEvaqH7SHL1S
sF/U9FGsn3I8YR+rkRVkFbeNKsivEFepyUS7lN+uFNaeY9QbI5TR00vyFBMImZOjAmF3aizuqUJm
XxNgts164Vml/nOUNScb+Fd001rlhfvHmQqGnLVD75HpxSp1l7StazK6lgYFFZZgoZh3zT7LOWPV
8zxvKYhAlNn8rUSj+Qf1jGX5ig+IeNbXymzTdOKQ91klTCp2un/mmtyq5zEYvmqv3HiXiaN55OCS
lFidaMpRcQUxPTSc3ph5p7Lm6KlR+k6RGvL395iSHfwc56SUP2rZh3meuJ05KFCQ2O4w8aowyjDk
hQfgEHvkOX9PCh1WZuC9+nvDdM/Iy/lOM9FmDqPMu+ecLoBaTq4GIg3r81j+iC8NcPfqPwXtXKtd
gCpkHWG+Z5LNICuYBmkkgQYR8UxKeF7Bou62A6yRXfUJ7xgVtdsLCNvBT+zw0Aa4LkcDm0DUQfpF
/s5FEIYC0tKOLsBlxZciKij9gHW9TXRUIR2oUlomMH8A8KT97FfFyHQlq5XvdhgjYr87DhkWBCDG
pkbLZ/OTSDypvxlIlD4vqfdobkKOO2AkEEGVKuYQpLoHvSegypcCnQiv7+c0LBF8Q4/w2MAvh+PM
OpkZ4pP9aMPIxbnHpn16xdp5MEdhoH4vsMhpwbDpdRk3zHGpoz65yrgBiXmAs96PypHOcPz5f1Fu
JNOfjyeXq6cFqIlIgJB6ftRBlY+6RbUxwYNTLLhqMBs5yu7m/9yj3K6sW+hBuggGHtQBfF5PyYO8
B1xkCeWOJD8PBf8Sncz6YlGwmDdKwq6BUVunGYVKEuq6iBYwShNK5VISfHLH3PFpbCQx9+dobrQs
z7S+UPI86+vQ1ZwfjB+7s5SroQbVBtag+jEs7l0ZlL9P9bC6zttBK9r+DphDc8NcXY0bIFJ1vJoK
12VcVAjoUG9R2heDB8XjOj+kOvXmbajnIaRVk8toKEfuP2D/YXp+7NC9fGUA1Put4ah3faqlO1eb
a9GSq8kE/zJAqjuAJy8HXGwfN439EGsLQoSky2bsxnOLo8eskkXfoe+3bs+6R0y82rHySM/amJNK
0GtPSBdV00+ZZxkDDd0BlaeAsL22cdlaYgnW893FteIi8ozDZ2VtmYfpfs34TbSZaC2OZeLfOAUp
vY9Kkv4B47NYylwadDUWhLyIHUwUiuUbQS5QBGMYf6GEVIeBrsTEqSxBZ6EopJPSTEOfxBot7sXg
oYRNcg9dJNlmFolR5E0TVJO2vPd8jw5H9k8zgBJS48y+PYHElxjGynXKz878214FVY7CqZvo2PvA
KCFAlTO6qBjbocJUhLMxMMolL+h0o6NV70qc4yPQP2/4ozu7HDmeQaZC5lvn3gge4PDfFr2cD5mW
twD8bZtMhLfOvXGl9BHAidS7v9sJUplNEUJ1XXjy0YvLxwHzkdsH5hv1XmQzRNPNhM0dRXXNG3JW
0kdayRjDktxheY7NcyQtltqNVoOLAkZTCluXcnwdGuN0P2sC0L+9xbTkrC99FsA5PWEWSfPFHkky
u64FFd99mc/rEtEvFOFtP58TyWo/WddbZ4PQUgmg2fqbytsBLAeBTZ3vuBGq0gTtkAZjNfJ8YmfX
D7D1n0DoJjtvlSj//LIRlti5/cwLoVMq86Gw3Ae6cwwMpJcBQ0CYOQPk5oG6oDdRzwQTWcaYPM9p
xmS+MhHmVeeWSRGTTIph74x/OjalP1q3EHf1uPd4nMxWsM1KKTbbUNt0wpml/TtNTUkqRPwtgoLe
Y5l4ls0iu8Y4j+9kO2ihw4cdmrl5+KzwJK19pl6+nhWciUfdtg4WZjVxYUzmWKgfTwF30AfClBOa
SaqVHXtRkurlGtvw3+QQQdpXL7W6mWrUr+4r4sgZo6BikUg/+tPtvSvBLeHKFqNWOQ+zb6ABmf9G
GLJ3YpJb14Sy48F2lrTwwo7PbmpEw8Nul47gXBZh0oId0f3Ncm0P56VEUb6pAa9yvPb/KySb1lw6
gZkKJfpWd/Pau7o2yqyCHM3BEkNLx6cnEEexYVlwpnxCZWZ0SMudwYreZyJDYHpSfGPbqusbCF/T
C2gU8RBtvgQWQC1FHGdkBPMJWhMA4i0EGn9CmegWXbzX1TRuOghjq4VFLjlj7m0fNBBr5271CxSD
SfYW2v7WDPO3kmDnhuzeFEueCw6bcg1sQgp3kHdJIplKFHyxDCYNFvwGjsk8qrD/vf2AOd135gWq
I+zIX9NqbN8nXsiL/qD+ljEli+Sc7MH9V7osyUZrWe94R/UM+RQs1JZod6sByfTLd3xh+wG13sas
tcoSJTFMF2pM2eVRsWap7dULPRirgAzfaYO5CQBh0dlI+SxNbPVpG+g7hhwOO6uFAg9B6F4mtKIo
MapWCmovrhYHWG5EyILyy2vTCdMeNZRCMFnNgdX9jDRU9AN1lI8DIcv87uiX239QKz7yeTD95drV
vZBY9bLktgvkh6HMiZEAfAWT/522GsoskQhDdozSjBkHAuigSDej9mVZrvd14WvdqxzlORR+9wqf
Xi7FPp2zeY8QW0xmK41wgwSliCTfCjolNu6F6FG3PvO5hxgG3tigIwLNQdDCWoD+P3GAmwHa3TAT
rxAMlCuvHloQc8hBMRClpUTPwAHZ1exnA1WI+53lho3knIKUQJIPpXcDW12A1G6FUaQxWznvImqg
9lhSCRe1SID2E94oSS4DlVC/bjU0eqtOMX8Z0GC8QuH4Fc2i4GCz1EhdX3hTny/2ayrQlByt3KP7
XdOreVXGr1fmtHrFbBsHp6frcB5mffVimnRZ9gZOED8RR6ZoBv/HsIZQWk2TG4jMs5vOhsowpic2
m5NE9OBn4nuiX4vM0bLafUXwnZtfay/Elyqk+SQcSLC8EULM3jGYaqc2ZOX390fSoVo7xwn54pX7
TLlc9ZEG9x4e6IRwdepPAjaWKLLTA4dILx7K/7rQfTQzQJpZEYlkI0yLch7E3ukqmG20zqmmLK6w
j+vIpsP9BDjUCRPepKuzWVHw6MVvgG9Nf1cUIJwbzLpJYzslv8YJmC8KvCeXIMhQKI480/Tpzzqp
0aSYjtJtSfgr0uQM7ne4wPYXjSv5QTxlQD4KYSJaFimQ1I9/e3BPX4oI1u2gc6GY1IqNKriflWs+
4YGDLb27fzeugPrkTtcbDKIzS3W0Kuvkr+Fte99+fLeM13RfwTf8lK69tFLGVW/U8gknX6fT/hNG
6oPHhJ1kpnFERWUHcseQEvI850WSF2rc1kMNKCUG2zP6e+6g93ZQsiYd9SyNuzVF3Jf1llOaJhwe
K2C06ci5selfxyUFAjotKInV5cj71nDIFzSOz5F7cKKE0Cx2IWyvKASUSo4WRM0q2wlY7TGu3idx
1adb2i5KKfDLV0w2ogd9cW6UAvO77L3HYNdidON0ctX+2moohCzYuI26SpMluc/y0lxvOq7x9eE3
dqPIQJ6Ufkq3KmBr6YYMCwHgB0RmA1+/a5nRsr0bBHiIuyw8tLUvpSlfFsJiCcfbma+WCcyk4lnr
cOcdZK9ZREiFk6juTc1D3HX3iUxC9ezy7aTJKvnBHLMdRCc9+SHLiB2FNTpCtImLgrTJFXYV/rhK
Ot3Mmn8XdqWC4xMV35LLAnS0mgACP6FHPS5R6I9w9PWdUBvk+qrImMp1jvXMcFvMMV3hQVes1Dah
q0cmrQohIK8kzHOvd6BYMgZPhVgj/pKz5hMKPq1JBDMKU8FY5PwvY7yCHjxvbdyJYo3jzSLsn8Gj
k19JF+wc9gykpUkagHBJMbgpp9mFKWJcH+ia7sdqtCm4d5pWMaJGSucCZ2P57b2KUgdchJOvhTYG
zMfL5tMqD+ue02IWTI3YuEXFQgA8qGPvOleFzL2z4P3YZqCUS+sFI8DdlksQcFXVhZrUSylBbah0
z37zL4/DXClyDEeBanKTCWvqTHt3NL4HSJ74IGUgWCqQ1PnUeEjOE6PCyflpSTucy9qtINp/K/1k
u3JNrSSYEr/1Y3PEesSvNV4DjVocsOGXhCugMndZ8lCEOaZXoLJZz8cLrY9vRFpudnL07eHh2/QB
6bqbVWJEe2j8i9IHKt4qpRwHdYpF//qWZ82uk8/Q4SedBgfFHVfKBc3x5HcN4tQQlXslzr1xwh8r
lA+dz10K7Fx3Mpq5bNEvpyJWDXdKHPiBy/dWGpYw6yW8VBcOzMLaMTBI3EFSifubzKZUl28vdkeY
pvtYDbKUzWEguN5GVMBTz4Qclldw5IYde+xuFAtxa0BvLYFrHpFd9S8u82WxGOpaBHAPOv2ZHMMv
R8yOzRIDlAEgLAp7oKxCFX/6RFa9yfgSoKzt+tO9Lz+rIYoMHSnb3RECorIOV60egg3VXcEppZ+9
qE3sz9PPHIGdOdZJL+qvHRLZ7ffRoMMXSNIOFUfQ4eHiKXQ7JvATlEXQ24L1+NRx1GQHDCOmBo/1
gJCn89gXkMNVKDuV3gAuQeJ3cL2tyI2d5R7rteS0qtAFO/zZNMASOA3ICcq0ZcyL1ScNElOQsee2
TJ+bqmEBTMX94eXZiP0dl2D7MXKpWbYp369KwEPCvzVD5GGk7FUykes3izCc8QRue8Nb5r4X8Y/p
TkJGcJsOGC9joBgE31UjwYy4K/etTrWpN6FJgS47CzGHsfQptuqYPR6JhpllNCUBNUS2K+DTjp9E
Gq8GpaVJB2EJCj4DqENj1Dqbht98MzT5BeHJ7h6Ktb37rVSBI970Ee5x7z+pepKJiFIf83io6wyQ
CMpc88nVBx9lor8ZPCQtQJihTp+u5C3cdl6xfOhceqLk131OmnlQrYMucfDVCCABrjpVIIV12Lzz
aHo/Y6/JAfNnBUlk/PFBTS58pQZ33l/vPZ1IKSpO8Kb9n9VaWAT2GfRT+EUs34spkORVRHU9B819
hesGjL6RcBVKeAaeWbXYw5tw3X3KZz7OSwXZDNiPSyloZNH/Fzv6yPS8/+uq7YPZKd0WF0SlC5gH
Rew750ws4y6YC/7VFTzqa0ep4hAOUTJ6zVFTtzQUoxajayS5el0YeEwIrjk5W6WNTECVtuYmUDRH
9hZN2+kqaa4G6t1XpdWiD30fZ4358sC86u5ftEjK/d59FwCX/xW/FD/NydJwn9rafhQbKnxHdLdO
0y+dPpc6s7jdC3uANfV/tDLwtd6BIFKTgkPfE0jH7MZft4lUXOEElKlDYjggYXH15k037B8ZuuLs
5Ft/as3gr7oRUwVo9S8Jeg+GbOxeFXRlI+KVzDydN7mQGl1a0QfhSFbYDOPWZoYbA41UgSENcGGh
uP6QQ74Jie282jTTj5UGyBH6KrYVIze02YAzngfjnckDEXrwQg0saVNrv0bEVWQ+uOtB4GLhxiAm
QAg16+JDkEkbsIu2QmrDWDt3pLXXT2T+IN3601obygA+aC+/+detgwfIJQRhNS4YYwUteKq++9FD
4kKJi/1owuUpkb/MuPlXDp9xDGSKrcFZOEhKgRxJWJQwzjsTcjU22ai4aKQpihOEEFRtG1POPeaA
NBsDDRQJ/t4p5yZvoKj1h8m4jpeY30HMkpnscqfNJfE4ok2+9gOTt0wSBlxHbwdNuig4KYjeJQnd
RHSFZHDCPQBdHlzUv2C2l0GebvYOev/LX832iP6BMx6Dtsmu2cQMdwp5Tv5gBYakIAwqwYo9R0mn
pcMSI0XoUtosCG0Cdx14LuOykREDrUuVytZp1ReTr08yBtaHhhl+4jiudc6EK9iWbQUcoz13skHc
ZTQZW5JRr3XB7UztETPv5mZfB/Kwy/UVWJgibZ5szG1Ky0RsgA+YOYTYiBBf1P3RQsUvwv3d6csM
M5pYS8TL2SSF7yRIXZTzF5o5UmDHIaLckYQ7cV/f8GyaIji3aFcGBmdARAtDHVQyCRq2hAe+B01v
tj1EYroqhgrwNGi4yTf6uWtdhj7zvytxyMCjFnVxqeao1AIXOwc2VzGKlVbuaWzAbK0jE8WcoFvg
d7z5+w86JR78PxOswTdve6LzD+GA1TBLkuNAgDvkzavxgQi1z9+ONCHGiDJ5bYaLQFL4Wt+YERN+
G2kVbuPsGfHJrXeJMdyf7yoN6mAKOHzJXBjQoJkrUzOLV+Mx8LN3Z81rh+jAxRpjiGVPD3LmkiKw
KXO1SA19ISUxRWT5UD5cfYwwVLOWXkAxMzhsTrXJLGHBPSJpDrqjFM4XPMHA46mQi1sNT9FcibR1
XB6AIIHKnsRHuIzjysLkzcUYy8oEV5h3B8tcAt58lUZSfXBMKNweCDZQRvA7p22jzV5CmyPskR/D
yygFjeIkd1onU2LdBIiJmcCpKlCNj+VtBXp0/yzuZL4vrlZuwlLZKJ+Aa7QjLHon5aYnzDtdLMWd
TJ+vaw9TfeZXwUtWEvi3ckrDYT4K2KO/RytR0LOSiVsriRZOq71KkKvcy/F+/YyVg8Qc1HMKk54x
8v990MVHG8ed19Z+YEwkplWq1P+AjTjMdnyVT/8IE3+KiVLpYKFxrler0GRKmBULeajcfJTi19DE
0MbHi1fJaM9bouclR+xpE71e4+wRSCQLC3B8UFWkxCNVp8IVJlxEtIkLsTexcx52jQ5cllCaHFdx
bARi4zhioJrM5CXhLQqZ5hCEBwVITRXYq95oxNG4195UcdH/WCmZD+XQ/dzkhPYFUqJx0bGFIYTJ
9McaW/sanuFimPSs6gpc6xjCbr3Z0cEzciaSTm3gpWeAo7EH4OuGkMxz6TSLcLOYWzq+0421Mmsz
wX+cYR7RTiGhFImV4EkW/T4sixUcadrKQKMA5Ge0d9hVcGzJopa4sYjpOiJJY30cEhdYGB0o7brE
DMhcPaFrvaJ5k9J2N8i9m0YdtgEM0mLSSZ1IZHF4sDFao7WzrdEQH/p5+zVxG03kxi7DOpbZ/2vQ
vDGPSzNQrGwB6Hp32KhZ/LJy0/hDvch6fB56buR+Spi+ziWHgGeO6jFG1ZEQhQhfs98wXSrHrAWl
1I5A1D9FzhROAFBU+53wdzhPrsAeBz/xw9ss0yfGK5Wn/4TUhbD50R8ZV1N/SiuhqJPST1k+Bh7O
PGyB0vVXwn2I05TokLtykC4kwOf1NBORUcqa8qvP7ggils8xydqqNBgA7JOcJ2yoh2MB3pseVQpz
CszzLZqKv1+a/akz44PJrEh9ehffpzao3odiEJqD7THTAovckG43Xar4MNFCprzEGmrAZdeKZSw1
koeBqiMy1EMq1ME++m9FlnHDDQq+brwTeoKJpJiuPJHnqijII5TOGzMazeNHx0NBKU/1DKgx+1vU
iKY7of6RJjeIbavypSRqv+nqEPR1/idvRE0ZtT0xiVyisPnLsY5q2B3Lv/YFAJt597vo66gZ6Ors
5iPsEbsnQ4Lt2r5tooM5SyWal2yQbyLtMdkXHJdHQUrmfjpfFqI4+wQsNkNW7UQ5PM5s8Hveb/58
8+5l2LFZSPGDybCxfFFa3L2dHsBkcy7eRT2UgmThSiIHsuCQUpicIXGhEE5Iy/wGCab/ux/uOIP0
fp8qnH1d7XkvBnKg9AsbPvTh2e/PP+XYQ+iPoX5Z0r8U5KcD2ImuguGpoE/jttnw2nC2i/82olem
UE0h5RThtBLd56/rCCAszQR2yltuhMlZx1pfVcAhaZ+stGd76iXnVAjbLOqmRyvdIQ9qxX9RkXq9
DQKTaf6yVYPbBdFrAbVYHAGVjaUyX0uscnLRnD5wzCYmpAMX7N58kDzXJw8SN1oYWnAM1/5fML3I
GTEZ39GG+EaxmwuCjyO1y20tHStDTTgfjoYWFjkgfSapowpZ1a3HQu2iZaP7uz6+f8T2+aAxsMZy
u1DuAKmnIEyTypZhdnsmj0xYzZ3UcVKZ+0/rdiRO/MWtJrXfasY6bRvBl3tnyLK361otHKdEKCLb
jBvTbMT9LyV5BXYy/yeT7kNQuCts45+rchZkp1dC4QhLpAqzabEHAO2DwT7C0toHXiNCWm+wLa/b
7BSjUdxRjaVRqoertX8ULNsySdBv+pMmfrElbxG81yDuxpkU2YGA5V+sZ+mtE/vfArX28quWysHD
tI9YfHsTgU2sOOt9AnABMC/s2wnY1+fKzypo76KQ5TgME61vDEQX6ixIbpSm7geczvYtQgM1gXzz
72s6rYzrOOlkUUfsRFTln61RwLM+OGzU5aF3q/4pcTrPmKW3axUQFQHhoi0pgFc+nHgbeta+3sM+
6zSGKnID6LCKlAbTH5MktGO0g3LICCeWyNi6AWGgVU4lqIVU+m+cRr7myQks3sojSiNLO3TMFIAm
Bt9ZISuhzI2167aEUrWogA0S4pd1/8px5rINbcIGoEANdDBvlbDNuL07c02HjMfNOKECuPfPx5d/
NPl8FnwGJwt+rQMdZ0SuOvfDt8o1CfNupL36BTAb7k/sk/gklZDDmMTCiTsSVE3cJb+5lt/RgMIP
2EqQXCcvCWYOI44AVCksLjMn0tsTP3saiKINksPZbJjHL4ok/y1xEtoA6Do80kFX/aXsHH5TCUJf
JIiUqc14LDC62htYShbnRjplmKDR8HIoA0ae1M1SY+YXtQm+B6r6itlQRn8n2MBF6a+sPfeHeA+C
j4bQ03rUR9eHMMmUvxFEBHe+gH/L1jLTxvwXa/XkFRsrKNo4UAWomkR0+l4y/Dkgu9J5npOMAL1X
t9MMuJHsixHUlCoVY0nKIhp0yuyYDVY6v3Llk1eXU+izk+OAL69pJDoan8ijAQue2nilvV2MNg2R
/f6+2+1UKkZO4HETL0v48pPMZPGK1QPR6XRPNwZB7UioSCZQtsWYaQW/Wif2pzhV/HLa8Olx6Ksi
5sJxD9by5Y7hVOWfa3zpcw7NMY4lkz3UrhbBGdzzJ7EifDUDoakuwEp3ILNbBGp35+hptWDlqoxx
/nlFR6CJ9NOaYtlrzIMAbOBex/xRpmnRKG8WtsUzoQN3ivH5saM0jRuLNE70nLI6ePdzgczRl6Mp
pfnMELp+MkT6Dylg4RMsKVZflI8PMOIi9OR8HUPFMbH8ztHj4aSvOfqR+QMoXreDJGIiwgWc+ZHy
CM9OfNMYdNm+2HKgX2uS4PeBOiKwpPcbYGLChYVo6F8oWuJX6BnOe3IxJOwC3tz28x43h4f4mMYG
vJwBz9A77YUcVT/qJs2BEWTcJafOW29BHZmP6bQ8sGBXnnb3ztFtnzo6o3gFKdJMO3ob+BZApppY
/aY9ZHJjSQRQu+IL0XJAZfIHGlFk2xAU63ZDkNqE0J9l4FnNXaFXIfjOXeWzFvU3pgRKgjLy4PP2
RvymbjS2VuWh6Sx39bQ10hY+D9IF0m03ekdYTtBgquqxqK6i3cgHGJ2tJmMOMEZSQASsTMkYZP4P
lq35jYbvyFhbwmMNvni5lg+d/nGyw9cRsKPLM7Q/0nDMqYw4y3pG/4ZsiXX3PdENqBUINd1TiNGK
l4ajBXt84V1Fx2lkw0X2aaMSTcjCiOhfwMv5DIPUDfaWe+ChDnEk51A/EdviEIgLm0kHbcRmD8Lh
Q02g6TkYHiLd06enAsGKj6mqTjfQ+deo6rXr7sgVVdKGoULL/fYxHcmsDWd/dEsO7HssKj8h+zpo
ei+Bn05+8qyvFXAEl5mu287zjMcxFz1oFeJlvoacZdl/qgkggwx9UkSAFX6Cy5FHSfvdw6zBskkl
fkjGF8pp9ZYScUA1N4kqQvhsugK5P9D9w91uRH2vJlbnOhsMm7MlO2yvUeY5Sqvfexdfeir2mDqG
2xT68tVpieTCqrrCmvUrSNtmFbPIT/tShR5QMQ2BRA3FWq7/KdIuETwhV9E4gNIM5+hxzmhi2xcb
Iz/EGWaDz14spnVFZ/oyj4D9YMQmsdSxfiql1E7v+2Vx2i6n0wTPhP3pFR1mAk3xDm/7f917QOES
r08xFvKyRylCtA2Ux7rcl7h/tnm+DR/3EZfNpkVml512TaFVSM2FG5WqfhVfRgFKOkj0HmvtdORq
ugBVAm7TQb1cdcIWttldxL72WUSV92PwTHeztzp1BB3C5/mF+6UUf9yDTH50JUXV7skYX/jdUx8T
y+4w+y/wSkwnp98DC+pmsnGOhqNsHXA2rfw+Hs19e3DmpNFCLpUPZdX4Tv6juOhBA7XvprXXuZo8
E1sOheylGRvRzxoviKvbG+dDT9SnQVbEtsnT/0+aUo00l+gKES1JyaqhnBev/ud2JcnPszP275cs
5T8gmyHrq+hfZnSDpIc03SkuL07X8CCd2x1a3GBZmPQkzpVxzmcJ0ZDbWUGErastQOYPJa3UBhnP
jRoL2M5R8rlY3ah+6IChpeSjEHV0LOMBU9NAaMoUCdcqYCZPgg/kCq11505Qpu5JBfx9nu+RGsLA
HJBrqpqIjTiP2D7eGWkF7PhXkqgGoVQ+oXMlYTRff4JItCebKUE+eJK+2OIF6hEJl2wNXhieicAP
1hZPMKAnlIdDBICwCCaGS204eizvT0keHc8Xi3k8vyymQMB6RlaWkOQDfF0/CMI4YMPRTOrvrw48
Zij3fYV8mcKTD9cuwvnQbW0yzLn9POpxB/fB/xgZYz+Yp5NxT7OueYX8irj3RCfzf1ss9Eu2CWfY
bWq+3kssvYolBHxBAWJkr/KDUgJPMzISvredKzR3yw262993rNigtHTyAB6/SkRqhrLNMeHPFVLT
1ngLC8I2kMvV6KCdpsofgrwMZhZWa8a8Kfc+qOR0g3huIEL6sqbM/T/YxSM4lf1Os2zu3q11Xi4S
ri2UNe2xHQ/MDZNNqi+YEonMKD0WanQoQ3AlKoFZ6HwEkUJg/AvTCfvMe4+uTQ+OA7DvWod9lLIc
jOLZRjMhF1GqR6Tip2evS90zFUTNLFk3IADJNtFq6Klfw4bOqoBWAt8kEAH+Xp8bvjjkchsR/oGT
Zo5nHNFjDUO61xXWWNqf88Hy2k96a1zCl92sBgDNm/8wEKvMqKGd6IgSf1IwoB6kMfZAT3l4tg6R
4SfiN/PpMuNfj/GClrOnGzTySbquk0qJlLKm3MR5NF+w8808L5VaMO4rIjC3p37qoTWI2aZ9LdA3
1Y5UecvdZRvDKGWTcuOKhfo+bzKASusJDCO2jkOGwpJRVMMp/2EMpDSSn1XuQ67K9T9s/vRDB2RT
OlWvvRMj35vzYHS97dsv099GbGE81MvjLbilh/Qt78ofK9rFu7WhFZPESDq/7qNfCf1qKr5I2GbE
yyW7Rw1HKBODHcG0C/HZzXd9dMAr91DWo4dS2yImO71PjEkxmeZ9TnhBuKKDHCW+vfdK7u7DhlbU
Buv3JnhEzLGq5ZmzSJNAkVYQ6bfqwSaQUe4xYgBM7lXGAgW3eEsZXbk6+0bMRcxRLFGqimA8vWis
ye15hkZvyiiXTX+2/ivXUZ4xEgRoDuKNX4P160GFGhhM4DKkP89+NrVyhuvV1EPQFYK0rokzl+ae
xI1hkWvdznLVstnPquGGgcXp2MKyhisqb4HCqy53yPl3Ufwg6pJ+01IiNiWh0QR2Eujv4MhkdvNE
vrbmRh+rUs0dwKizmgyMTZUUT/x1d7sDVOEWZS25rpJASz+7AwvbfHNhtj/LakloR7aXQthP2YHU
kPJTQ8DMdTIfZja/USXc1zV3XmW/TYhtTFhyjvVF3n7WWF6Boi8EJNOrZOE4DqYlXMGCZ1AichEI
7A5AkNZDmk/o8r72PNSW6F1Um5MYUu2a4G4IPeqDYjpBBb7goQC6/X7hnuWQ/jy3fJtzK8nXRI1c
hAC5FbeOy4qYLhPEaOvStHBgVeWC43U7JLHxhcJLL4f3FkC3HU70ZGKHoKGa765eMOtIDhH+7P1M
d7rTNCeK/KuUoKrWgbs+DjVODN+Pix2W2AZPdjU2o2aZVBkAnwAHzwHsXu8W/OTRZGE8i34OmtPq
0wQETtsiwPGsdVln8FJtatJP5B7U5WTN3F/RRwmrJutykPoD5kkUgHgcEOOb2GFxoqn8vglXRaSR
WRgn/65//HVwbdkvNoTkrIOJOLHYfz2CridNmGeItopMfSrbqQvZvCCIz/BS6Oz/huRd2BrTXj7C
avrsmzZOQz1DrZN7nfP2oaWwTX8J/pbHX+cglNk1eUouXjy0VgY2a5pEOzEnRz4daLxRGSP7rq5W
bADaIwwoap/CL77moOKTkN1wuqQOiQUcVOSCLjjdroGmxmlMwrTZ7T9XV+ppV86ZLCMEMl7yieGI
R+WMn9eXbckqGx3zKlxmfaOJWgGgJdcDTXZuKrJQwAcwpBgY3+DKPMejxWj7yOYnKCCtdOtRaIF8
NG0O0Lf4gZ/5IL8MfyQ+gnpUZzADRb2b4FOqsGyXe9Qcms/AsCIJa61uT86JHlYPOy3XkUxw0mAF
n4ARaJwkkS++zqNmtcUolEakmW0pjxgMrrf5gCyn2BkpsqtZ1nZZwdsqlmHRXG0NxeDreVAQLyNW
mmn3vLij5AbI8rz4uJ7PxlfLuEkVvJl3f0n5H+mhr1/FuQyDKnrW5GGpjKj3P0Lv+bG5KRhaLO+b
7P8JIX2nVPtFqvIXJgicGm2Tv4K2LgDZzIqqEjzglozywaiKrpsdH6K4WADXmwa4nuf0ScglkOkK
BD25VYMkVKaUo7osorv4kOPawr6PYv795LFbSrwaozIuNNEtbJsVX6H0aSyJ7uOK5zfxARFKpSEy
fvDDvwP6rJIBNuPp7mWUNYGOQstzMIm3Ev8NvyWJytB9Tr7vreXvxbeeco78dW2jPHtYVU2XcYAw
6M6EzkgdiMykO7bZB9f3i28A6/FslSBPDLrUU0LEN89Ih8YyydnCYJGHGGTJfD9tIrMDklSV1q8j
sehYwlhC2utjRqpXzJpbFZ9JBW5onJinEIMM365Y+S2ozibzgX3l90bkrKU1AvQ/NeAd/Yy6pDck
laqEgJ6JreOaJXKJOwAmDAaNlieLEbX+ycnKGXEVPILDA5YeIc51s5e/YH5b5VM+2y2JCy91ohkv
GYL2an1wgaXUrgW+AvH85+bNgjF60s+Qfpe82V0wNpWdliSLNqkvlpDBjW7374PGGAGcGnOwB9m1
+ooXOA9svIvqTDEOS9yELSZ8KD1Jmmlt7I7PQpMSvUlNm6imHDuHZFgkoxrt/HGOtrZ4YOq1+VPf
KbYdCSM/Sq/UB09FhWDWVFwyxLTQveGnq3Y5bccO0zA/ucXqNqLbmEPBTnaB63MS2XWC89buYAYj
L8hWKNsKppm0iY0xxxRhO1mtkgcuMgLoJRKAO4S5Y6KKRLmLbN6lTLW37OpvWKYYVjguanqj06Ur
OiYEw952kMmv0psokVDXh8bTxgq2LNco8kv24w4pK0aSFPMGaLCZC0r8JGvpmEvcaE9JF0WxsYOF
iWbT6X36e3T4QwjeianrKayKFvsCrbQ7bIyw9L7CT4EN3Gk+NDX2lHXdVHLtZbT38lbgcGFpSU8z
5ve8kASrsL/gaRfjI36lIdys+pQ0bs6+mSCHW2+9ad8nmCf+18saj9R+C2q0jzPoXetqrwnm2y1B
ISCMWdcjFAgeQDYS7dd7fHae/J0Jjt+JALjIWFoHlB30ofWXZ/7csQQEIKZQaAAy1pAwfP/OI4PS
YfWBDzk7xAiqLi44D3QCRMLagLt+rfZPucPHVZv0RDt+fn1jjPEKhFXA2fuG0m7xMF1Emejb6MrO
XENFb8z3YNV8ti5kzIEYKxXmPq7dTbDcZLDLIsVaW5svOw+P6df/aTGfRgrIQU4MAssrCHcp6L5i
KW2KNz/axH6K/HNO6BKws8OLbOEJQ04e0AimqQS+PpEOjyGW334c+C/6VUHNrKC/ykAEMXaV978T
/d8eUEjBwnp8FlTYCmts2NQKpeGZy6W/rI1rWtx2CZoCfXd3FPZyM7HRvBRnaVZX0gc2MBYm1+lO
nMMq22rDyIBZeEgaHVuE4nzAYsaQz6FNUEDxNJmbj98IQxojEWj9WafrzbSjc9fXSZ+kccH6NoqA
t0bX39McXfnj0pId1r2lCXoxkHjCA76+LNxwkzQJjkQ47DYJWRIZTLBN0Ir3HI4N+769WDb8Iwe2
beD8aCSfPyeHLTDorOTIbmf4ORSWeMhLvm5+TiyyWAZfQW3yK6dAsuzTPEhlZLqq8UDYANlk3K1l
mCMDbVbN12J+bGBtYx1FTGR1y97EvtGklG9m3XQ5UqFIhhgZVj1njUnnN67qfDlVWlHABejHTamC
Pludh+i3J8r16XiBdwaQcn/Kqd6cDfl+rHxoOdWq8QnjtWOx6qAgu3A0NUKZKCYVwLcpcGFCvDK2
mmolSMC8oEp/LSwJqs0zix6bCjS8ywdRvfJ0HnTIPpexwnfCRRDxtRL0QU0BSRUhM5jisSsKoSk0
5QHBGmoAuxOMMcU2ZaKJNfSphG9KFjlcHYwa7U9FQRCnxSKo7H/7lDW9uZ+fSmksePsqhGfK8HpS
qXlgpgkVDsN7IT3XdKuJK6f03BTIMtoNoYRrLCqi8g2bd9eXd+tgbkelgRN/tAo6Ec6HDHwOrf+z
hi0Rw3IXJgb8Fv/q/tTfluRNdvf9ubSqYL14uNt+dCeaUloEha3SPeySerbZGyktUrLl7Cybx+9t
8f/GMBr5+7JZR4mki1QFVqb1S5mf+tSLSeP2AZUZEnEGGVZAF/E4GFtxE1S8nGWRiz55gnyncVKI
7VHPvzfIG0m2ipilOKdJVOSRq6Mr9ipF4tuE3mLKYtTKsptWtOkEu5U7rkHv3TV3OIcncU9YYkhH
aWLAtHgv4WgUmg3DlC7GNmss85af0DaSA+o4UKiRe+7oDfR7tGcPumQ26x8yBz3+nsh9mRKBKZy9
BBseAXVDB9x/E/6cFzbKuu5kzcd2Moe+591KSGE3W/3QU4IyvkUW8gpNifMp6xumeTkFNMOEjLZn
KzK11K0E9DCy9uaWUhSURmi9rb8AAvuVI2gKV/JipwKcC+CL8NK2hUxz6WRbXFU5mANtvxmlrV0t
FFeFMJ+afKuyUDwUOqVN7a137AZ2GJb1a8x0c+sqEiqQX+9zbbzkxjO7eIpHCiJZNEp5Ai6DUDx2
9Qwx9aZ5AgNTDY3Fx1yA94MhqOxKviBn/In7ojrjsFQecsk2vK2DKMG6v4yMrmnzlvd2RL1GE17l
YIYFXYajg+HhUEieD+PbdHsSzQ9bAvKJEzRZlwk3mNiY9uiNrpkyNGAewEmhddzzsLXtYaJISFVQ
wbTros0QYmpvVv4+T0XUj+TznOM2kBkQXYq6TnGeYEW7co6/i7IOJZoeLrk7/OL260A3X5ZkSP2o
/FqR1lZmYGU4gQnaN/3evfbXQ+bF9TAkcVEjHg3etg9F7PpYFPbJX3uZRQrYDxe9qU+32c3qc9cE
ttOijFbKh3y/yEcw0xHjxzjd7MW817vmgoeIU9+3o+DrOwvJDj81BUJ3bqxW620L/3O94TELC4mX
UYG6Ewgcmh+aa2mUnuokBU3HRPyEraWmnyAYJdXPSV8We7HqiWBZu26Hin8M4d1jKkhCWGV89BrV
JNiwrEwqr5HFhMjUwusIHlH9SJzmcefj/FNSqYlhTKpPkiZtPCF6xkJZCbUUUVLKM3LLb+rmxq8r
je2nt9kz+tbtTpCaUVdvMmPl3Qz5f8pUp+ORN3kQB0ThkaR+mU9Jfh8HAX/1/CmDSV8h+LioPWLE
YGld09CwNj95ZADMIW1kcbyeV0LV+X1jRbdLI8TJOlCw/8SqLEtXJJnUmixH27wX76mZjAwzagq6
Hfkxg/78JLvbSDoLew5a4joQPydttuueC2oovtIv+LGuIcccSg96i6qmbjRrbQ/2AynS4OjdLFoE
85ruKfZzrfy2v6ezc/6J7ZVpFxZk39242tuPmVRBNz+VOpVA37kQr9Ypy5vUdy1gtDUdppUI9FOn
1Uv7YXA+ItGcnldUD+nh9EQAG0tAIT7snFldvf0tYou10xGlrBm2iV4vY08PsP35CdTnhQiheoda
BVBbxO+D0AD9QEJJ5ezuWuvJY/DXNGZZJD/DuMISe1c9uFqR0BhPTuuYdqsi04sd35tsJNLkBeep
do0rcorYdVa8eBi65hpiziekV+1WPNx9Y0HgpTtLJO6UZPyuEU8ZXaJ92LjBknEvjZrTd431UC2s
FlVmoHdS0W8ZfOuCyfClbHZFEV/9ylCqi5Z/5s8RgasDLGmWLqGxrgFSlHiqjIREhYyTh8GjcJdp
EKSJ0q8F7j8GrCXBCubnccyb8A8G2uDky+XWoWacarMTYJP2+W2fl45WyjU+sT9pPKo01E3mynMl
XpWYKnxo8J8Bxg8SDA1To3odl9Yz6W0TWFxm+hpndJT0abuwoZR5cHcwn0BSRd1zg1KT2jHzBKt4
q2AtTCoYr3l+aGk4Xgg+dAOpIUaGOlxTUNtvKGaacjcMatEVuJWaYNRp6AUitVxz3A9KYjovwFNb
Aul+rHjHtFlA0TI6yX3iBwEa3bFB2OWDuQwBiLYE4M5oLWzhFtT9At8riOHl81sHbkupvgUOD7cU
asUb97MnvrlNUMfv7/rwmMEAWBWSbq9MEFLPnNqqWyFXcXz6E7XsV9UxeIrr51EdLMlRQdlCHUua
JeYLlTzMgNO9eN1NYrDg1FJLzEHeDJCFNGL5YoH1zqIjineOTeSnbguHxGexV2xcAzU+zjt2JPGd
rtZJzSSsh5PrrBgN+ueR1bM9hz4SNV+JGjL37Djz14CtwOWbxbvB1V3FGPslJ/W2Q+9QKs28yKgK
f4EoiGlm46swYnWIzwnIFRKvehyekpJ1jaOq+WZfqMutNORz9HlDaSIIovdtLHv6RNbFQqh1sfXD
EJcCbmxCJVNlWGYSpSXZqXwG/DEuPaChA4KwvnkkTYrQJKIXg9p/DqiYpcXHAIbFTvTRkoc8E5SR
kykrtAbSQ9QniYXK5moHhHaIQSkXMiHXffuSzTRd8+KierGQ6NBJ7A7AjTaCF8HwE5Xiq9UybTXR
oW3sN287vg6HWuuFgit1nrNJRFVtor/oB62iXv38KhUPw59OVRopedOkWE69x3z48+7cyfQij4Fo
YY6wNVNBGSp23XoGep5rNodFPXUihCoooWXNIqmMWvKM7oA/wVMAzj4Gduw6EgllAL4qzawroMrp
gGj1OwlGoKCmWDXJzEGPi3Y9QjO5CXQf29c1PxBJMtgnYXzWOOC8TbCdp0RrAS0NyTW1Slc77Zg3
gQLWZM/2PnqlZTJHv4BohstEGCzA3nf9619leFxO4yIvzjfA0KZIoUcz485YTijKvcEuQOeDOtp9
6/Xm8IdpMa5oDEnFnXDW93FcpO2Aa50ayXhEcVMJQhw0C4Nqp11Wz9GJS/ecqkRRav+sTF/WzMW/
ZqpGdjYxxyJXp2URVJ5MMGdDWHnphSAz4pNiQ8g/x1VsAAluLBsj4Yqt0QxCbjWBvQRiQxtTawcG
giVw1m6P8thgy4ODcUNf7Ero6z9oVPWoWv5eWI8bq+FcEgqm6e2c3IBJXfcOkXqzesH7FJePmrt9
jP3FR3J1MrCChrOD6wwu9sMKkRoZrp18e/59D8GP7A5HTQUYnDna9aCGhiBwJ2rRNOEGYOYKkxPI
2MVVMBgaCv4vSqGioZDsfIjFQD1iclqEUPYTik1hnPjCzxTTYuYXb1/TNxOsVnCwDBYOJIZRDYzD
MfVETdFzrKXDcj/FDnJUxcl3bkrb0Lk4rlyVP/0fQslpg7u5mfzgr3AREeL17K8I+jTzEQZPSeC6
YD2SLcdKIkyG5iaJ5aZ6N9JfCTBlvnhrFbOd0ut/UTL3rORoaOdDN3caG6KJuXg3/bYGbkGZywwL
4teZrRYUyqgz4/my8H/OtVISf+KaYrYTJ5ECar07NKuwFha0MyjUCyVJMazsSOU0rUd2iUcT51Qr
iERLwgKPxEWXnUeyu4JV6HMKp33N3eGnuBc1Y6Q3BZ5Ca2TWRAUphdVuycNgsGHDvaG7PepDJUiC
5LNX9iAIlWFOTlGcR1HFnW/AULU31ztRIFu0yWUbdm6RZS2rO2DmB5ROcLBOHk4eXDkFYfk6sqJT
UQMBaB89VmoQGbIdnbSTtFpVdMPeZSYQixAHX47XP2LCVkj8AI+fbCVJDGdifCjbi6k/0ZcRg7N7
zyPjsV/S4ug5qK6IuUNDXfZc8HKhKJd5RIhBW8RBsOS0oiA4QNISW1Z8GGzZNqu9SnkFPDszzdnW
EwZE6RUmsmKi0FTaIMcSI3jRCWpi3Q1ASA1DVQL3RRbFvgiowpKrRrOHcGKsi5xX6puh3LG0sbQP
ZDGqZKzypBFtxRIxzzRZ+eaXeqV0OitYwO534G4fLN1pmDO4VSzj0aq/OuWiOF+dioGERVOgEcHw
OmyIsPgDKF3l+NY6gMnVqaLcWNDhs9gGFBcFoBi22QfONwV7Y0ZthwKSD3yXoo43LUBKRA3IYjE2
UCbm6jPFYIgfe8nyS6NVz5mo3Li/a4lInzs6WOJO7y+D2kqQHAHhbQ5H1jmMMFxkGnL+fOtwB+4Y
X2uDFVSkO0uC+kwUrR7YiyKAmThlVbqFuLL4G2/2xY6P1LXOFSaikzgiJL79CVa+BEnUWubx09ZO
J1rGTQxf6jAnMUL1d26jgyvHI2O+rsh8JpcrcfXyNw4Hwor6NiVYgxWlRnTVq358PSfr4Gjun/5+
+HTS2dGOay5+gDc7rppRB7pBQQMaZkDHI+lYl1v++rMH1tXDUgG+C8BeY+UIFpFpSdbXHuOttdL3
f5GbD0p5ns6vtnRU3N5ZwfY2tlCLEkw7kJ1pMorfGPIDONUMEXPwn72/rt4NyjN6NGOpm2PWdF0D
p0u9LZqGCw5b/wjghQIBLgSvOyRw0PpYtPYYW+0T8+SBF49Svg98A49PvQfgKnZDTPhOnvG1fwhm
uXfjlfLDfNfKtFYy0dos2N92aHsz71mhhiie5Bfe6uZ/WDfDjj2yn6fc7bjpXxgS5gONrywL0Nya
YmsGg4snzmuqrRCT4BFXeZHuekKH9Ft2JqIPn9z+fK9sM2/h/oUNDpIpe00PJTPeFID0EIrXye1M
4iHLZ2z6CypchgihRVxxD4Vy47QF6SJLfBb6T/EOrH8du5+rDO7V/n6PrKoWldBsYieYv71fTxPO
93tzKlQOop5D9yYKrlSgJkT2JSQ/fkElvw3HQs+UVmMrrVXMaJzT0eua3pvVMRVQP7w071EaNUZi
0KKZJwrBEwAjp3xNmzPA7llsGUjkb45C2Ky5aMfrr7BBwLoKPNDCsLDLtGs9bprlaxDys0Ija2bh
Br6ywFago/aViZrfjup3IAeY7fx5ogI/k4zlmgovdRMDcul/HjvJnkX8zWhVnGnbMicF3VETrfdW
XOHU5HyXQBhAzttGg8OPLCOA1UAWcb2fBfQSPHQlLlv4Y1ytbKHAXC75zG+Z/4JfFsCAKhuG/6MS
LiWeT3ftYKpDSOzJ/TWIp80pAtZJNImuVQJyylpdfMBz1XFyUo74/VTi6i/eVWriEvbtxBE5+HDU
p+qnEVaVTl6VYWNBHRx0+xHWfaqBcHVFKPCDYF+JvYTAgdWikhqMI5z2Fen0mpvN2a41FwwIkb7y
qYixbcWA13hYiGoLL2MSosbPQUSjTeQtnwwXz1ubN0F7usbPHERnlF8KBCgs1ap+TStbthKIGbr1
FwnewJI3Taqxpa1OGZGNBxki1mfyTzJYK3l8zP1t4yqVHxSYL/nAfkUkAocVEFRnNn5zIlnE7XaJ
gM2HYxnekZgWtJvvndl+ExKjRJs2lI5tmgwL1Ffdwkf7RSnU5+XWyxO65VH9RMHKTuIh95LE/bsG
hY/sSj2WimKdck2BAD5rVYiDSFAmb7XFP8AZl6TNpi44OA2X85rElkV/cTQQ8CMju2QoTe+zMa4N
V1hU7Ojnd0zQZ8Y684YQ1PyMzr8jCjKjJwgN5DepoecIKN6P7fQVuV6QtKqHBoUZIf5AJw6kElzY
Q6Hq9JV3M4XJcowEUY51q5Zn7mHZp3n4gB7XXD5N4fRrlihpSU9+YAMLdCxFvHhETZbr6Hp0cHOE
DPA/msXc0jy4QzmicE+c6alFkkkbVorsMi/aLLqDeg/1Fdpb+YRKi1ZDEbfwMWMcN6rrI6UEu2ES
YEJrLXu9GvSwgdqXkzHxf6A7zajQIPtlx45oorRTu7zaeBix2yQ4klmfjWUXwXFCRiSJOZ1yHtE0
dlNzQ1EfmVQ9a0iyWqU/fdpmedzTo0ZpmPW0asB3dZR7Ahs/WVCAdIIuxnyWpAjA2oohtz6cAG3F
snNCZ5nzsqGkuEiLp4I8SeuHbnex68/sXcT7QKX1dwBwc7nnBm3MwB2wj1K4L3A3khSCP6rxujy4
78yeFzpb56S85Fgiasc87+RWkXjTHr2bLQV5zgpnUcoQjbLTZ7/1u2fVOMjvLgIko+BvcgucX3E3
9gEH3tbgyxg+O9dOvfnP6qBBX5QBb4JlXSeMemvghbYGevgX//HeB0UtMcQD2QpJJVsDRoLOkJGe
ATI/p9ZaelwoXqMXoCfo3Mg6rywwkOiJ83W1XzF4CoOFs69+Gz9ybqAy5ZYaW6EMTMwuvZ/U5oSl
SORoPSPLvkaDBYyNJ2E7BtUVZYtGtFUT82X7j01u0ix+MAMd9DbmyOLnpCq+hgTamGpH80hdcYQn
447NvmUCSVh4N/gkGArnBAfprPJg9J3MtgkOsT0hnhIiFNGhTZktBgrqO6kWTCF9GKMxIs2MSfs7
sx0O+Q++5MKH83bNF1R31zhyY1RkqnrKa3dDNNrffInvj+8KL3GKZm7iusJNptJ+814KWtLoBfGZ
NNOEZkZ7BVU3s26n86zGrybgpx0vHwA4eeiNuOlWHdOCuHZf4iF71dd0pHw8jL6yaG5fVN2pOZLw
6Bo3HbZ0niF6TeTQCcSRwIcRrKSIheSnQhmiE7Qzr//AgGFzHbxHlR4riGo/WkGseDgDngVFeiKk
KllQq6DCcbB6Z/FvWE60mpdRNPPUdyz1GeEGViYBjIGF/G/nCZ3GSfnhAtUkhT+u9/LVfI01aYZI
1mq8P1vYP3KVzgw10qHS4YSwCl+ysASiA6exYtNHV4wKDiITL8+RQHMzlHa82hUAa6cAo4LVQMo+
udY77lVzNfZcT2KTcwA6XiKvUVoQNmyyxQQ8EIREvgnqg7NtSob9gCzzWB8P8GKMif6V6SOL4+Oc
Zja/xU8tLCcpkoIwC1ayhmJA4YfZqcfX8lu95fN3wvpUE/bq+GGkPcN9+mGGF02s78dShYQkbwMy
hLC0rawUZEgWZuvNi2QIQeGD7mr04GYtyxm6n1RODa73tgYeF9hub6VlHrScnH3K5ia8jJ+GzAuY
pVIJALCVWquPIw5vWcGK/JCyMn6mgZDNRGHSYaaLyBnJbTGSca7jfMlL17t0JyVGb/upop9NX/Ke
tIoZQRjOnj4dNpltL17kxPwRPFoxCZf0FkVXS7yt+RzglhZYBWUQv+Uvj9YzsOkiniPhxbJWEGRD
ueerqA8B0Z/cw2jN/QVIelFkxlTkC+l3mc2c7qd+NLUcJMjfI9Y9g/KqKsnXaWW11pFqNFXAy79x
+f7pZU3NSpW7PeBBELpmnUpHlIn4logTBmH2pDQoGgySwrmb1FLfprkZrJ+BTH3XxOeEXOLWNeOc
NYnL6irA57zmDFQIwyBlX5eie97z/Tb2jmGrUuxu1tFOIuNvUbMqgEm3KTSLKuX6IoVstXjO57I7
YWwb//YbOcNsVWcXb2PDY2b/JNIs0iEuYOsHaX930edEa37iAicnpVNLb6V1LDbwOlmGtwqJkTbp
qYiR/XG+W1YpeCFSAt6W1/72sdLDY7WFHWAPTNyeDXDkiYJVFwi3QzcsBwgflFwbR1YMdXIaxB86
fxyPAv5W5I+9CCb66HtMB3U9Dld971xKTgbxRNbwAxQfxyW+ahbCTTblU4qgl+xr/f5i3DfBaS8M
A5A9olj0REQ1faW186NkRL/MBZ97fauLy2HLmW3HRQcWF3IVAC/H7o7mUge0zRgEaS1IZAy/ztY4
YB5VRKFcm+HnvqX6JHkpsSLqNhvZjmFRIJZEqQ00ZF5iiA6rJdRGhbqh8TeoTxaWSPbr5l7G7qIR
Tri8LR5SfiXVaboinWrkFB5Y1az0VD+wNhn/27o6UMF6mkShYLX/MjTbp6OI6ZMqI3Ll6a7pCJGc
lx1U9X7mNoFAD0smi1UH8uF/ubRkz3jK2F8VnpgKaBBbNmQOpe1/Z33Df1ef05UaK6HeYIom/wD3
s3k0DubsKACcqKKRjtrC726RSScwraIsKCBVtuatoZQj50aKs0qjSeuK1gTBrcjEo9RpNt8nQpob
FzdQZmox2+qJSbS8qNU2BbueRKjQiaeRb8b0TzAxEvcLlejfPW5XrH+ZVewYWto5mAP5EbWDfLYD
y7WIvr5WDc1RqsLhVdhtNRi4nTeie9/baDcyyuIvVhsycc0BvkXk/ecquIgA5MIDvV08CdnPJ2Dm
BukO2bTY94r7gDHwhfH+nKMFro9DxBZ5hnqXrkSu9ohHVAtiyoUL8cYHpp8MMn/uyV08F3NkLARw
XcdG9mZKvV3RHErrNK2smdFeQFUUztwnwqONZE6L14I2xKBAzKuEDZYs3jsI1/AEOitlMHRv5uKr
rLhNwijHEwOz1/sdgbPMCfOupczlkP/slZfupid8jhPzDaf0nqySRn+y/cBX/irIcINR16xRnEiC
OXWc8JMboqvm6XYhjKFuLmby7PGFHyDzLB6ZnUpOvK0x2bDsvIcpKH9TmWoqU2nXCg9PvVwtjkNO
OulTDVT8UsuAawJpGPSsBhERJPBZog2jNHUZFgifYIKMtwDgdTyf+v1PPf+dr3OmCxXQ8jV9e6cx
DLwpqAOBYaPe4u0A1OrqWjeq4cKHVBimOAWZZUc1v17sMAGgKp6Bmzwf+zE3larO4ARdEe7HPnRQ
lHYYdRDdN8QX2+PVHMNsblb7pDXxsAyvtEIxvVSCN8MwC5aUacedX0Ud1roXzdXKd2K1q9PS7ref
itcHXAFU8yzQyHYd/vjGd75emef5uOO/QSY9FeAL2mPk7V+Yi8T4odlFZLnMSm5h6VwAiJqP4/zL
mj+aawGmfOMzAVMvSsByv5K4kqRY2GlWnkaJipaf+tiZnsoJ6Q7LW0HDdCWiszPfVge9tsehL7/q
+G32O6nh5OGjLSjjVuOwfOTCHHDAW1JyYjs07bDK5klTXiYdR5qxCCtMvBbk2Yn/RZeXTkciWMsI
4Uo24XGZYrEkUzG/FThninLZUSFlKfWbY0MAryJXshAUCLZCKE1LbXhvZt4d4JBOsIyRsEelTTDu
YPuI3vtGhYS4SChjmgFACPGYHhoO6w0tfkfsrPpwWFv9ISGmv8twsgJtzIBuJ9YdfQd4xuxNYx3f
bzeqI/WRrWrt2ImIV7mV0t323foOozdPaVm5PDKnuP1ahN7O4pjRDFD3yevHco21A355mvaSODNw
4cRyQKzR8M+4C4XpRU3Xhwhbdm1+nv1Kq0n+mLsfz9QlXMJWEfZPGEKS77LxMjIYq+Zx8yjpY9UQ
IRSrabwMZWGW3Eu2LrdIqkyA76sVUZ1rPwALqUN5fycZpN4yGBX9U/vPFZeGtDUf0A3jXNHtzFE/
3gO8X1j7s1IYyQsBj5bS61Q64TP8q5EyxQvpwMLFVzfsZ/5XSggvtyVHrboqrD0EufRZsxyo+ffX
yx+shpqztNn94Os3AeS8rayrXHrgEenk9S9aeFFcqyAL35/824uG+VMajXOeF43JjW0sj6+gXHlw
WLivn7yIdChRhRFGrr6poRrWL5942JhzV2H86KmjgTKGrc6kEfwFxppeEEtcx36vWAixmU84LTxD
nkK5s0dtyQPAEdWHE8SVjtmjBZA84smpUjfCsCC/fbElW3aYuWZJlw/3kaZ8GlI0NnJiyhcS0ZyM
MojMLyMwdbLZM+FywnME7xUWOD/mEA41Tal1FAYDGWGSgDndAcYKwJe0XXjRCb49jK6YsQ+iWcen
qIFWpKrIvEtGDUcxoqQnjarjmyYmPJSlli6R0OhSaWviJxpHj0q9J+8oXALnddPPmXHoZNT5/1BT
3w7q/Aus+T7hDxJ1wQtDTSI1MSwNX+PsQV/Ng8+H7OP6vGO25Bky5veA7TD3XJG9e4WpE1CBg0u/
OTX1JivxjPouae3MIrKID/07aWBcMOZQyV04aN/9PUtzWTgjgsjDbc9ih17fVjfuuAJOCxPESbNf
Im9WhadaSEqtJyIMQbGp+Wf4yKl2dp687Ylw82966hCHA4xC3FCNbHUcsMXy+2kWD5R/k2Vq2UoT
cr/H2FKIFvSw6PK9gWSyMFECUW/7WsxDisFwnBgnVAOITCDZhd4tBlHEZeINl62iLxuP01b7Bs1t
sXaNBdMxV3Cl4JA2wauP5siSjMy+Mq9urV9xs3EEkzC79FrtLnVQEcyIYH9QaXX34UJI61QCYxA9
jTXc/lh0/3fIHILaG2IxKIDHsrfkddskuzQHniXbvDYucAgkQhlkiI1nIIf9/nboe5LslG8LWHDU
eJ+i9MRYceIfGatHQ7/85mgNLZ23rEIREvBYHMWIKdOvnkOoYuUseORobwVcviLXk4uy7iTNkp6k
ZH7+YmhXuCsrLt7QCbP2IASgZwHGjokbsMOP/fnfgUFSqqqurPFBXFPt8kKChxQdoy0GmxDrZgQx
yFvM/Kx44XJiFOx5Z6fjlCk1IHemqYWult8pGmm0L0PU1oWxQ0FmeoeJHwEPBI/lpWmiarsOEGuh
h0BrrAgGnYIlPqXmrAZ/OKpTtGnSflxWHObqD9y6L8yLSgiNEd+jPst/V2UimnOqRuDy6y4SN3ei
Zw4uyFDr4TkgvjT3qgZqTf2aIhX8zE+fs6D2bfLbQPNixAqjqq7ydFA31UQpKlqQ7ONsoJVq9LZo
48VlLOo7mtDRyG+Wq9w73oyDt/qyHpTLyo/pS03Js25B88v1b9fqcTmTfY+oCncpU5+ZgvODpvaW
FCEN17icLnTCoOkZkjQJ6n4zBcWHCK2usVRaLtjaoFnRT/wwfNz5/JMnT3Iq14vYL5K31pqjVNpp
9qnYNNl/zs5TpAALGxFlwYiYRAq+xK3tRUgX1Ixdp0n5iqspXfmsA6UgwakYw4ZNiIPjtqbXj1Ut
xLGZyEahWZk4KfJwEB/2MR8w7LyIR8/KMBsg2Y+AUmpj3A/HBW3ZamUcc2aPM1aaon4tZQyt9O39
CoWSR79HRLiLzNkoTOkaVrqWRG7pYpjql6VEulqf/DZdI7MTjKT1YzL5e0aFlXrCoh2vizhmkaG3
P7ztLk0+knev5ib+ZVaVhtQmGbn1xoDgUd60o7UUJvlRIjFclYUB6ZCdL8UC3oZ4R30ODiy0mYc8
Ynf2CQ0Ls1X9IhV9DM9Z8iC8WuELxdOj/zkvxO4VLqMLrMF+25l//jvNquOtStoMmj+RcK2HnmZa
ZZzacRzTxXMy7mW4zGGMbN/vuhHPTN34lz20MpKL6yEGGHRzsHUi01QOfAAKhzS1Yjbyh3FoGuXh
M1fffpG0ShL2wIcKLwoaRgOEOYMUuWQS2GW9o/SkeZUOTB09SK7EEYV7EUDG7ekVCvoiFaCq+8us
tLYWQOTCm5u4eaGtqAinINWKI5iUgKfAVSRTiaPro3bfIMElNcpmVhfyqkV5Ou6I75tP2qLPmBA8
VEsm6ptXftiL5mT+FcsdgPcCXsJMbKeMAUtjWgvu4Hn6Fhb/jESP2vgRcYpFsks23Z9kZkrqzn5x
6ssznQmN0hw2ny1v2KcHyccS9LatViOuuLRPVATPMDvx9qL4ITyM5i2DX2uYo/lKDuKnJoWznr5q
O0Cfvumz0yG+dCcTjTb46SMAMTek+W6YyVN7SSLO5AH/LiT5ET5yTmhpk1aw206lTBY6vR76rucB
r+jQf1/WKJwUWyUKE+znRVT8vp6IvP5NYn6wrWL3jZ1kReuZ0usbYwQ3YCS7TEI5QB90qb1Maz5p
pSunZpuzbHeWdgiT8HpwqZbtJ2JOK5hFgq9OFuvznPTc4S2TEN0Eq9NTvg16bwMS1VDMMFAa3sMf
pwEaJoztvtZZRmBEWgVvsjIZ08uBv0hNqIcMwdRpAKugqeXhgMrVsXU/c4Rb0SOarIuMWEMh0U3e
S6jvXDE6olzPFZxoWpq7GUK3nzCPPN6/wtIYLHXX5GvuDbfRTgkymBBsn7Gy0yZxqSvb8Th0WJf3
deXu7wC9CvUUBm6PyWGody6d1k4FvFQqEZ7TFamEz+lSl9mfkyECfC/ixzlXQ/ykNwhfB5MouT2U
McfsYui2ujuB1nS0Cx1VA8e+SsMlb/MxQDsWBm0VTr7Y/GUvzxrsNbBWI7VFwCyMraieBm1btqmU
G+tBwO/fFz5XhuhWFSOj5b/7ulyCus9npw0ck/S4lWcvbH1tbu5SgQyIRXgthu4Tk4fdwRNfOajP
p03vDBX/kC6HV18kEcU2H8kotlKNk20BKJ896QuOzr7Ig4o1qNnAKYYciNpvlRTZJMh0EqXOgahe
E936w/oEMVTr1G0hSafeGvWtD6s4UkD4sv20m/7uFVOy5XZvfF8LN3XEtaJGKcMTZodQqWvAf6WE
CUP/Rq1kOO1qQrT60qBKCbhlpG3auD/IF76JDNTQjuOfIc260gBBEOByXepXHSu9o9L8MV5i2hJZ
XHu9QyRy/Y84tf3gWisS6Njnx4w0uW3tEE/VhGj+0af6zFCrq/ZcRHOlBTbRX8s61pHQJzMuQLK5
oHVttYnwWMVuUgkfuKQX3A9EhsknbU+Xt7cYnjn96MKxLpQj/0gbMD0/I3UG4mYcxU0q+wkNTYh5
fwm7Xzto4X7byYkKL3Ba6dUQarvHMACEJ8l28opbhkP4kDq6I7A1ECHovOQyJp1ymupPFw7UeskK
1i+JU4j9CLTuAm6ngVvWOSDDZESDOe+xAQU2Bs8neVb2PhgAL4Sy64yrtgjcoGzlEaFuc9IoTewr
bnI2QLf/Lzm9+auF9axAFLeZ27YhIrq1g+3odBFggT5vz3u+iLGNRb6InCbSVHlNiSGZ1rkbyiEb
RG/AdJISDFKEOAre73IiU/BMfhdlCW7gQa+ffP8nAKQKbzrpdhNn/Osr9NLfF3uDFezlr/HlU0q/
0N2U2JnTQQCZC6pZPCFSQS38RowGwijuAYmxD5BxfQJLa7bowUPgV2t4oR5FlGbkAdMIVvy2JbTM
KIjXp4RCWhoKOjzHYvUWRZYfQuWfb2SZgkdlirZfjxOUTsJ6v/Mku9AXbBRz6UVanMP5oSVXq502
SVu4/oz/craF0ANK1P/AupB/gV05bkR3XF3n3VTlZrYQClwKfunuIVKiNMzv0a+9g/L88uTQ+YUq
lXwb2XL/UYKIwE8XfP1fANv5CZhqZnqN5qm+R4wmVPwKnB2c1gxVY+4X+oxQ/rE5qp+Z5FKul5tG
ss/1UdnNc8OS2XfQkGgeU90PdNJPZq8DWIurEcdM03UJCCMSQMvIaS4cY+UtyfBc6c1o3Yqzukz2
J8f0UX2ZRX2EKc1nSEiLCGqO5Sx4OBxfgdIL7HoB2HZzvL6x7RqLnTVvgDP4uopMs4asXDw1WZDl
9UFw0EHbkChoPO75Wv/Z0Qdn7SqvrhBP6qEjVD/gJJv9fwgOG3cV3b7eQVAsqxXHUqpXx41zkyUT
wyPBWByWSMIrIX1lpQt+KF0hKb+noK2OP5I2IIa5/ZrZOqPfUWoiAjbnbCPn67zzEJ/solonYn/K
NevGak17UZD0a62KyS1RsLhVMWfD9Kq07lur3O4vPolxaGOy0pIfKdKXKAprCK67CCtsIE2iHU7p
+Y/lynl74NzURBfktWBN9tvrvURlme/SOyFlnfrDxXdCq9N884qLDrB7BSndAkoTJ+v6def7jPLk
mqh1r05pZmJ588DoIBxJhAeLXvun/tjg7MgG148+OSCEZdfAZhbAhgHmpr45eo2ApUznDsvDe13+
OMeKtXSUg/omq1xsqK4ELaKdioE2Ee7d3CC1f/giUCA1uZ4L7osPGH9FxxwmNsQwK4lx5svAX2SA
n7zXLPyxfma7AtML7AfHXtXGC4UXvqRcuXUq97k3J/0inX4tpeZ9PC9E9chCp7rJVTmAnkcC+PIG
SUI9qmdLIX3+124wF+9HdTDTvrG8pFsexbmHVEtP6D5B2RDKCNFLJguekbgI8ACIlsUZ0yBA9YKp
HPT+IELB0T+Lb9QIrxRpeuk+BgKgY4DoH/lNoHMuRAUTYATLc12fcSmpf6QjOqt9kGhuv8tKYzHY
Gw8Silh06DXvOWiJPZLVeoi1/hOwmgrVz4SjedVB99Djgjq14yerqv8SErk/dw/gb0ofVd87aSqi
xXYrWcZJ2O27+CYgOZHXI3T1CNx1PCksZF5TtjPxeRS/scKbVxShtbvxvPp33eIVPzt/gBoJTZBO
x2qUxPEM2CSDRfdhrP0mWn0gJXYmjfdGrbOzqTthBJCTiipGoa0KCYXJdwnaUtUcKtnhB0b65HZe
F/rRBkuc1gZZfTcj8qL1kBMBYRapr814ZWFrkfKqgYzp8cQWo9XQAzISpzwcoPaTGalN7oLtwiV0
yZUc2VQAgFsqiirdw+5wDXOm7XSjawmTyPC+QQbtNTjLdjBQBN5lRMurQQRGx+JTA+Snm1XB8tRu
tiv1YLSFGkhh54vfaVStqkvlQKLYg6xrOBH9iqugemhNjDqLHGYPl/YhMeF8g2yS1OQSsVv2b66c
EmLC/nLL0GOhXjrb7mbanSW9qHUOyIZP3z50t7fNwOFJR+d41ZrMWweY3v9Zz6BIMC8K6x8aA8ED
n1FTn46HJn2eHuvjRAjSSE5MzIT/F3p4rYI1aXAq/MzoxMRsFVuT7pIZw8CQyl12JKbZxt09D4Bv
pa5lMdfZXhilL8dyOvD2NQSo0DAOtzorZ7OsUpQvKiN+ASgdEUQ09MgxwHp57zpczkxNf+ef5qtp
bLlqqOPgncuNewjkhxBTYFmIRsDtrbAq0YQUkqSUIAmFUHM/BU7YUdVfX19eUSpjtf5Dyv+LetQ1
dlkubcjtWI+/rQtMMT47KZvCH0+scD/aPvez7MxIs0PuaT439OtgGkO00qTDkm7SK3g+IUuS/qIA
8qeeUVOIbn7YJ4Ov5xUgXpFURNIvtJhsHWUpXi/wGjvNZZGg2Riv5d/QirU40890lKN8sMHTKeov
NDTqBqAGB+m3stt/2lIMX0KI4sP+vR+XRyPQwmVRycJ1YxcjZdna+LkiatpKjh6AXh502CrrMImD
AWDQCcPcOgDpihx2vTfh9YlDVt6CjbQ/WDvtXNN3SM4O6TRY9pZt5TVFxCpAA93JHpKPYWLB8Bxe
8Vjx8M6fclrWMDLNgWrCJmYcnqkGfjCNavf3TAhxf6a7jbu5OMJ5yvWeLHNLTQ7ruc9N9zYqvXIH
+RXJUuCJNLDXvqYfZ/Ip0IjGzdruptiwm3uwCMfXixy+CqgrvquV2oLY1DpGlhx2Ooi/yhwXEMaN
DhCVkXIMwpXqlo3L9cM7HN1zPjxge/F2c/GizpVsg/9bWs/9wU0qqCtEisTnzS+CBFaEpgcHmP3/
6KZttRpC+rULqfpTN7X1knLDg8cQv6rwRCIrRkFVOFZx9LEaf91uR/iPFEoxaIWgjHSEB55flt3V
3ONyfWRSCqzzP6h4rh6xYNavGKAcZyLWPtdeFWeBBVk3gFv/vXuFvc86dTZCfV57iaf5gahuoah7
kUY7KrXNF8us9hbb2wEB6OrynDcqHTrKE6wAhnsPaaBibS3BMJW8MfFLz4nRJQk+pHwCGF4d3//a
PxOZeHh8UOsqKYerCY2c0dMs/Hq++9TWRlAHPEqWUkg0plipUjVQbXw6pn0Pq1XocosIRFeXIXMY
9EqvRo5sPPnIgJsK4jHpqmUEbLO0Cdne2atPbrF3yayz896XHIfA/d77GcyTfKF9PwBtlWBoUUVt
jAa2ewBTMFefbEXVj89UpPTAXC93doVdVCkeBvNFOqkiy43nwPbQZSjROshWGh78d9ELdl6BXrpm
6SlmlNo8ucd4mM2IH77kjbXj2dVlkPBfZnaQ6da94E17YMbLUOh1YVPzDczUvXjLv2lgZYu+uB2d
ryC3TwMYfVAeUugPCU6eWfK7XdUPKTjTy7hbH82avkxpwTTaQUydY8J6vMTFGm8xyLtBVlrqUzpa
P91iIZ+VtzShrv0ysy8ewr4mQKzi6pX+rYyPOlNraAg57sQgr5TnoR2H5NEvpJ6p+GKILgFa/fWv
ViSs8F9K/6UwMrDthpqIOR4bjT5CPv4PsMMX90hdaPf67uo9w2VudpbI7HptzsulmMnrm9ywLaKV
K3n7l4yv+Ldv2+aHJlOLkuRU0F+nOLNL3Wvl7/iYumgmUtzFHleXqOmsdGd5Mvvxmc7QMoi63lBQ
2ljm7t2NqgfRgX5h1G42aMECKyF8y7P2E+DwVudGXpYHtv3qeG7KVjzKhfEfEZMnZD4C2f7LAJnf
hcOm/aMmbg0TBEPTXlnKZF21tPEphAmUFIbApP4FYxlbNG72xNusPKue7m20S2KdDZq0OdkuFxx5
1MkNs3ZCjrWwZyjX/3y01axqEThdyr+66ooAe0cCwv0+UKM+/tZM29N54qQaMlgWOIHw4PuO7WuS
OXTx9GITF1DQASpo+tizUKDncd/hgIVR9c+pMmErNkMGe0Kk+iNAUUVQ1w33sbv9hUHzF/AMvBso
6MZ+AfG2HfS3HbG3lf1MgGAUF8ib7eK+EhoBtVeJLJ1CnRJ/6hhSCJBjYCiiy7ot+pI4QgwkeqGS
6QGLEcZWQe00FNgof8Cd/TFInyA1VmGLmUUf6kk9R7LQ0L26BCO1fxjRk25bNhDH9/5I25uOGrej
a9P47Y6AYbBmUyuSDzcffFDmd0R3CEDhtHQ7mqRVKzxdIK4ajsFF5qS+HlOWCDnkeCUyK+s7gUDy
lDBIwfRSN414nbLw0b6Zc84fSqBDQRJHiYZVo1GPfkBudNcTXtjb0J96dO3KhGUVAiT2Up88Aq4U
iwAfcbEPQoKpPWC7wySj3PDmdXeXluclLPecZKfJhpHP+fpmwP2Vw2XeJhbMe6T1Pz6FD8E8A8Ji
D0xcz3FICR5amna+FALuU37FP9wpZr+h0r1/CgKUUJWDfT3gWRi3kqtgsWwZP3hsnu9VkF5TivuX
6BE70uHayIaEa4ZbEkdtFG0TtJg8PYKpJ3/MKKx3KmU/GXbrUn/0BVvVO6mXQLeHTxQr/A0Yvcrk
cJHV1xX8HD22Wa0Fc/mLFUPC/jGUU1cf6/0mpRYT1z4c2tbFdVd2aVE5lb5uTxSX8e+IrZdprgQ4
Veqoi+EVh8YfwjhMZGYYDCjb9DNGv9mcdIVWgzWa7nYY/UOKt3XZibkwazBnG5sMdorCoCem9UF8
3ndXlBkQzvufchtDAC2dIKvaJbqxz1gH/ACvMzsQDwwCxtFA4nh/aCloo4ILvLmLBuHhJ0gRZpKL
iW+/QVCx8ZcLLKMkCT8oI4uMSNySLFBukaHv0Vwk+BakgQSqYm3g+uKnni1oqyzB36tyAbhCNG6t
4wv31mI4qytm/l1sm6cJA2/qumL3F/naDTUtwQUTDrKRLI5SnGYC5TUMjBsl3EvcwlULkivvbG/Q
f55tj3nffgdYndBN8xxcHUgy8scYh6r1OHrFmLLi1C6+mXKzt95MUbt31+yMs5oM0w4gME2qF3yB
awAWdHyfISkhZllQywkoaaztyfcsmZ2LKeuOhZJsZe7YYguXH9uwxKKpFMrA+EoN05hxMvmRjg/M
eeg0qA5aAjg+RftqVTQ/JWeyEg42OcPFs/1hqPkE/QakAdbL2dvKCRsQcRX1XRIbkLwiGpQa85yC
aGt58Z3G6xFgzIDS4ZZdCHHEE3AszR94V1r3vTM6AX/ELwWEe9kQPBgYNnqKseUAaWUQVbSC03s9
l3F1yFy29pCdiyY6B4B+58+kYVuJvJ1ik7S52InR17MzyqsDsN/N5ily1myVRCgk6UDA/OeWbq0L
eY1CPY/Ef6vKt5MEIPuTFthJ8eNfFeU/Q1/3fX2xBadY9VGDVwviTKKaUD2rdYrTMbnEzqaaboht
19Eu+p07tmWr8hxUIb+FWOyzMr/64LmiAUTUprltabjFgDI3cC2ldOIsHJDUOod9jvTny16vgus8
RPqrRMSK0BJdB6yPWE/Jc0Iq11Wo9DpHix+pwmsoNiQnZLl9aCm0Lu+5gYJcIDAYw8WsGBNGlJwr
q/fkLkbteH5DsSKKLqZDK+YvgbXTi2IlHqWBBwdwUryiwi7vvKqYYa9frrYGeuoWA++KzR5keOet
BRskrKufzGWdPIjkljqKMkie22RWsyYhC/ahZLrY/r8mR5AbvlAjUPql5DJ3Y/riExNaRUtUtdWu
0HEsCm2HtowrVmkkfhwjiaZcilXXGuDVbh4HxYSdb1boffvaqYodCBPGxXjdW64iMgznsnwLY/r1
RhpaGtDNBgktOIpC1J7p8BbyY8mQtBMj18ihsr8QD+VcK9Mkl9q4TEy38cXkoNIhp2gvUzxYyJec
Y1yJfuYlPygwia1Op3sOwJ5w5c4+/0FI8Rd6kAdxp+X9HuceWmqS5so53OVY70Pdfbws/JXB7Ryn
h4iB2uEGBqDhfVww5oMPI3yQimyrfuQCO3Z55f6jI9dvSGm/4UDDe1B2DD/kXjAqQP1Xqx3hNEVm
NmqZZOnqaTmVoVT17LKQkFvr5SKiT1E/4gnoB7aXTiqQbB1Bj4wOpk5+WxGwA9eswo7bCqB/YACw
RT0TOu/PeDgozktHelxvzkfghvDWfn8B8xZeCGeExOoeScGY/NBbXBpEyyJm7C8jQVs/N7RbCVVy
hRIMpMMdl5K3DgcWgIuZcJuiGZnb0NCsMVMMCgH9TjsvtEs+N8cI6bnItPjOicXCJAUc+kyE8Qso
6qsiibqmCRCy8ORH9ymeJ9+20PoU/bzqnqP5d8h9+Uw9Rl6Qr6UQ0RWBt85SFBLipnwkaR4zjCfA
iKXD/AphV49a2opzzAOXPXZCskYfYRHv8ev72mnoHJdgEHelclXfedWB3MjMkCMYVvL/i12l7AM2
OEhckxgl5f3Ut4keaT0oKkecKYL5gJWEHu1/I8mzfKaycQIWpGAwR5SQk3Y7bIDYyg176AmIkijY
O3mto4rQyYj/sLIJ4U9/E3F814CNwxr+F6vivl/4TARxACnw3ee8CVxkP3pM6q3U5VLNqlb4rBjx
dVVNz74tySuMC0hHOHps+6G7Bn7rMT2tIFJzT+5uPSV1OUNRT/nQJaE15b52aLDgRr4THrVDSEnZ
vLJimdqY8piaSksFSiRbmvJqZrNJpWn8QUGbu32URfjNwvD2v2f/gDDI08L0spBmfhpiSt/tGQEX
PVktTPdM9N5lEH9MIcYoNWPXjTS2PaOJE6JO9R51HWzPoL6sFG9BP17lVyn9uZ9zhV+Pln3yFHo7
deM2rm+RMW+iJIpVKnexjUBRwMDtWTQ2jYQLBDH3wIwqgiSp7jQ1ShpBeFP2+iq/LOU7nK2aXebj
ha8VhT5c+FSxpA54Qp0m8dUsi3tW1TiezJm7txR5do/YASyhbwWle7MLbTGIAN60m3r+NmBcq/r4
WjAwrw/n2vGaZS32jHDjn0yN3cMzbIxPeTAoW7b9TtLklLRhqKJqAMhEyVwIj9RpVgo5ECmwPidG
rXJkcaAEJZZPt7J37XMA5n1ykHdnWBtCSbYUf7DdWRd2LxXISyOnqiZI7/c8aOQmjOv02vMy64gE
zgmZk0f1GR3Lum32xHRK00rG2c0jtBx08k8vd/orwxWN8EjWi/8HfYZP3aZHQAqWvr8YhH/dzwwZ
oAXW8HeGRMmZC/UqnlJsImr1Qlw87dPfP13E7U3Qnh4fyhxFKo34SueMKTMJBg3gvIXaTxdDISL8
fKp/HG0XdGgTMpkmXDqgWf4qwlt3U3ZmU+CKoegf98Y8e95Vd6tNN2JEZoUWrPP9/GO93KhyPPMz
LS5dCmyG7/bFyE7MFdXLg02OBVRtq59YvHHEf4JFhQPXceDXUJfZ75NlEHSpkFiEHD8zpVBfo+Ip
C2VYbNaasQzSCrobET6PMeb+XTOkj8FGt39sysgq+rpaqSa4Naw182t5bA2WJ8Go4idJ0co2jM7N
fNks++HQkZWf9ipi1vxz0s9hUVCH54pvv38DVKd4RlIMJwZhWw0L6cW57GAcQYqXwGjT7iRqJz+S
JiGbIpM5UrGG+N79x0Z6on2s8UEhNRzq9H/GUfzenv8/HBCt6/cBq4qTZHNQkhuFtQdgCKQwnD++
uB+mAV+dELeEJiNcP9How19xBCOHRzr4FVLX9N6hyrEsYFdbzwkk3RLO5EKKlXOm4gcIRRX06Lye
eN8OhxbvXfv6jE+DnhxF+Ac5H+dUPuxFlTZcETgen6rSL2o6JFBFvbYDK3+FFOOEzPJExLiZYNVa
dMJhbmHJT4HPQ8S92Z28gS3NfaUj1LdwM5st/xGZeGnSL1ZDgIHcJcD1bbniwmPTrJ9yXORJk97f
960e1ALT9mJlEf4Sqhs6762ugukfpiUtCGnp9IVxQ4j1nLUPKyrbpO1QBZOnTV1AyfWAMHYviNB3
ZJObDCjT9K6sZIjBT1RazNVV/RCYKSKG4JBBxb7jUfp6wMGAAhyKWLusC/ISqbucL6rP+SR33TIo
eb/aE8sS7mUSfAuqwdgMpESlBJP+Gfkjl47EuNiJvD5rqNjaqqFPF5PfgtaOL24QDYzAGZCzrWba
p+rYd349w61hIV0Hvgw7CTlmd4Ta18L7/et97uyw6T9nOQsVQLepns8scv9v39sR/5BZ+zR3wAC2
t4mLh92Fp2ZXQgOqweyIozRao5ko7Dade5kcNGJOxboMtLhL3TNt9f85X5U9MypUotyom6SNL+A9
jji1JwY/PTxvgzsK8o1nVY/e03EizELT29Xk6EwuMDPAG06vYH4Rc4hKi4MjvIlN/tmpgBfwuxBS
O8Qeh1yVHfL3HEfbXm7AOQ27M/6C8rlXOSZrCQGJwMPw+cSaSfKVmklCaj1WndIfdTCuZSWwuOw2
GZ0BjAma8u9Ij9Yugus7pTDdcEWkbKKXAwxiPanLG4h2sga9+Q5vTaHEDEyumdtVTw283aQ4yhnL
qEk33tu9dVDPi18w8c9lKCfHy3PyrHxcXz6SWPM1HArQr06TFyaHj3YC8iO92PaEY1znw7VTiIcB
2Yt8RSChHAFqGt6za/c8priRDy4xEYTfA0ses4hAfwYF8wpE6RPGhT2szK4ptWgDoDGaJ21AjWTb
+ZW2TMv3y5oVZ2Iq4HvR3j1jN6HYM8uiKzQOpXKDPWGhDA1yfkq/w+H+VnsYOqWqruilk9/JXA3P
Q5M6WGnW4p/wU526zIHG2jqg4Ck2I9Vlr6TD/hnXBl+Ni2TIBQPcDadwCf8u/ZZPtCS5/e36i3eO
XjgaFFSlQc/DeKzQPGz/OfDzAKO59RXujlHFRxWT1iqKpbNABYwwezvnJt7t0vNpZDZJ1kemZvbt
PzAXgxVe0EN8ZiEu2JP66c7O2cLdTIurRa9LwFoEAZvMtCGW+x0k+A5AK3LJ784gqcIitvsqq8VG
BOczs8FWeGaSe/aG12W4nHSWoakaOJ2nWoxBlId4h8kedxuYu1uqLZtC19UNWsQGNhIwkkGeVYKL
+mdKZOfwxETv50yVDJl6jvrsm85X+yp+xmN5GTaiWN0pUEu2pEiop1u+uRlS9IQSUZU8i3SkkyWj
cb03OadQ0M9lHzwfaTAHICXjpzt66Hrxay4v031jyd6CThQzCm2aFCWhj0gFOum1aXmLfeh5RjBU
TS6T0rvemuDV3Jn+ACPkxfz+NKeel83xJdekz0spZRKm/4/PLiPGXSKo09KCm/TkV+jUZ+PTsR0u
eZr4BKlItLE17ihSkyY4EnQzrR7aIUZr69sdza4qfXLYsaFTWO4LT7voOCl09S2mkeb0Etz4EQrg
Bxc+c8zRVeMKBxtbMuqhhjTwG2izAuujY1HWdEi5fq/aIlkio7rK4H0Yvh959VsKILopzwy1Nc5s
CMoh+EtPDAufFJIug8Xy5WDrgv+9qGNJ9BTsHygMFAjLo5M2tXuqKBDTsf1thj8y8JQmya/2tmTT
Xyp9clh98aE9jCcUTZoJL3phlEFFSbmH//k7kLpYTaUgYUBsoNd2bJSU7cASGiWR9IyadctVgcbL
g8QY266ovg5P+AfzQ4NkNl36vCCTMDUJMPFZ0vSvRqiMIz30lawjbsuxoiF6lh+iKXm6pKnfmbny
KCtHZjHuPwNQKKFJmFyWxGZ5hiy8/OexyfiDpbsYIpyrhyeCKcK6/g4iX5rKw2Rtra34Tn2DTiOV
NCdPn+IvQuGgDXcFeDdrjxi2kICJarZwRHbSz8WRdfbIQN9+p9hbCEySh9/4YAXxBdwa2q2EAnkg
K0Ho4zAUi2jNoMy/fFQ6v+HTW0TIZrSOvjyfXDxcZ4UwALR3xGvs7ePrVo3wL1c73MJCp6SW8/z2
StoNS7pI75+qe67lQ6kwe9NwRNtya99KnBWE4J90S52DO0GQYrmXnbOwW3dwc7tfQC+rK7+VGCfJ
Jj0RyOc0dGfBbYh/vyRv+k8Y9oKqQgog4AbnHUTZhvn4InbGr+aDP+iH4E2Da73G26UkKc0An5ES
Wj6MAUmW9X3frEuDFH7JRP0l4+J/JvCI4AcALCS7/JWJvaS0iBeUOriPKY4DJH22PYzlfhCgoTDx
AixVg9uVdQH2TZaZra8mxlLz/fuL9GP6rzbXvj7NDqXGJuGMM+0XIGQLjiHI6nPn20j+KCYDas28
oZpWgpfQL4TCOMvFWhmsWWdqhFKlzSW7EsWiFB8vxgeO17SD6oo+2ySRuLSsXsD7e5M8Zy6ZmvYk
3K2omxJKSY9HlB63YeAXesvKEgoAyGBG0/my+2bfHLhZiRcg4bnxsqdLvl/NtdzcuypTpvShEIi9
CKxJ+ppUzFUfxIHaaY1I1tWWSQNEbbWASU1yP3JUe3+o3zckceOdlOu1sCfIgxWOrZbN9IXt8yeN
zwcIzeaKteP2YfhQHkTSA8fLRofrBrpW36Igfv3JkXwmuX+BZl45SDySPHEyXEL2gwODCXpEhrjH
lQ7i9SUdIqUGaynYPvvBylO722qOT+ttOm6yQNWclsNmf41gStnd4pdcJ1C7vlp6atxHruvgXV1N
NjfLLlN5qCEDU621y+R7UjEIrmDOYz3FgrH/AywBe0yGx7lUqkgMkdmdI2gDZ2009vcF/D03R5FV
AutS7cGIDI75+jIkCXo6OpSdd3MEdjaZslm9qCc1BD2vUe9uiRh5iA6dCEwwh/IT3sqRh9C/qY2K
m2myf7INGYPPtrTV421n1FovFogerNE0OGpSJxiq7kEzTJfCHE9VIJXI4w1GC+8xXdvg+3MQuF6F
ZsSmsh9HZFhyGS0pmUmO5SdFTC8jVn3goN43dOdPrq1K7LdOSqN87GCA4G9RhYoBVKF7z/bciZ47
9kv/dvYaw0MklmeuxEwtFUSiZbVVYIbUzfdU+MPdBsNoZfgV5zE3PBGuoIBzDHBb+ac8uuCJpZp4
jHqlZ398Cjw/mKXGRWvqF5C7P8vZLtIIUo74Fk46Bgu+8DDZ0MK6qguOqPjMg9hZMnQIJdJr9mJa
yzcDqvxHQU3TqSDCR/+4XalkyGlE4yESd1gqTIrrYFnyo973Lolf99/ChmhLS41g6LmaEpVv+6gK
5kc8P343EgLEpKrAV6S1FibCK4GigFLCObNEymkcsqbsBJLWtrs0JinS4B1eaEf8Pp/+PFDtWWtD
4jWXqqFzkbfdRzXjg6rCkT9DvkKJ0bKZJok6sMcxoEa3Dg2FeOYORGElPTpPoRTMZBhNCdwbVGXb
Db97jyPbN67udQDt0Jo6IhuzMdWyFW/P3VFWBSjOemDCQRzB6ScQqd+zYGls/gbknBVtxOk/g2u5
kPOTS1oCirBAGXwMesfHSnCw99X+RNRzy9Dptsp8NJkM/YBVJv0rbeZ6ya4YNrHDyLESiyVioObW
SnVGo2S0FgEsLuwE7CoZy1ZThiCxtp25AM/2rNrdiCfArtySozn0dNEyIWqP121sTzkyxwu40bi8
iTgHtCJQXZt1m8HoZqPDvkJKYA/rewz+sjK2V7YZM62BFY4S9ey3qAeFNWPCpl8wqbUMq8BF0GG0
9j7GUjKzLNdlKvvCRVLdZ5e1REHwNDOAdZhEZu4Hn3IXBcyUvVJZ9/mg5liwnMs1MSreEIh0uif0
Ken+66F12g/ram+HhWKnCJrDK6zmsPVrE/XmW7JF3wFcmk3zT4/8XM1CoeYudV71vY3EUknNBGcn
vFUo4dHfcwP+FvC6hhrxmwND02QkbPIbaI9JQCBPyRL+UmAB3tQdLtMdPAIGojNortycjppCG3/z
df+CSUE86hwbWrRrIocQ/wAAQmDYh/4jTxKFwUowBq3Qxv8PM5khwWiFg96RU9LWTiYoCqjPHIfd
vPOzGQvUFiE0jn1esayhQmoBH5wAfBRjkOcx2QtCpTOWQx+oij344ezijnQRhlVIhVDIfrvLSt1K
CahfSOLnuQmypVFsFPjoO4FCqsQD5y8UVL8wLuP6rB1irV7z9bV1j8BvxFgbfANDsX+XZbSHBNjq
YHFCAGvdl1YThnK8JWh4YT84VqXovZf12lXZY4raznVcP3E9WmC0FLBhYpog0Tv9vA9JjTMr8cHo
b9uj4jFMOtS6H/wwIslxHSCxBKqQX95OQkytrrJbTaArFLUo28NVraORASjxE9A4eOatKHWfQrno
BR6yd+ykWNLr3TQHx4x4ngw3FnM+aAipbScwAlWTxmQIjKxGy4K6lI02pTM8OEkQ0ukpE+yRQ9ZM
CbgJTn5n3jedFdKfn2l73eBOj+YpR0XDxb5QE4p3SBUXBUXE8wEdo+4Pth4tPSb3SrgeE9j9pFjt
G8T0XUcBfBkhlzaOzSAi58HLMnYBOfu1zsZRoicguGyL30UukPLRDLXrye4ScEA5alku8nA/3zml
xR/Oljfsu4FHxX7oGWIcpqj0erG61tz6oHJ+HcBY8DtryiBnej217O4jRXBxenOGGT4gzbUDqaTV
Y+GUZFHNSDHlOmTLfBgrdxPTIV+wBl9YR/ZFgm2aC/KC0bZ0QGPlJ3oXJXv115XsbuDQxB5JWABl
rdFsknQ3HslXN3Hazuv+9loxqYQhg/lJeKkHS4XjwyH8HN9hstL53y/UFV7fomipp2QZoUnoaJUI
dIRpC0HyaZTdZU4jAL9DRgeCpfA5Slke8OsZqoPHrJ3xs2Zqd4SDy2C5XTbh7O5/mWl6X/lu1WBk
Cs5cLIZIqpUCdsI7/jwKhuND7VmF1MoCZu4kP3BuYi4qfJyqQqSsrGH/UIVm85yS+iDyDFeV9QZM
fxtJvabnPFDjjHPIobHgcx9kpx2Bb9CZTJnvEozvW0GwY3OOTWhnH5r9IhzP4DdVaGSE+kSH/UU4
JPAsSJceRyN9lBBLWEHitCz7J+5y2AYZ/G/jjzcpeTcJHyX+bM08udP6WoPgOwWKfsKzAJa3WdaF
5q+E8gaof0yP7ExaLXmc9laun/3jUILdsD1GsvF8OxggIr7m4eUylTNEQRARbj/fQ6tUT4L67Rns
Eh2M49pJGlzUb5u2R+06hNvXBh+eJ1H4GSgyBRaPHT95VaSxsx5ZHlk2a1aNHo4TlZR0qvmJqBou
HYxslv4C2/Dw82B34j1Ltx46UzdedcHIOnOgdqx8w2Yr3Lb5/oeoYEoFLXHMvW/qgQ3KfvVRhpEn
XpPDB88Bm6sCYbBSEcjED0Z32fXgbjCgEscq20LL3nP5kcEIwU1CPORYK5UAmyJZv/nNOhrIq26k
mvs+D8PtG9ShairkAMoo//beq+iW7pH2E4ZJa7V4xjSCtjElIiaYxp1GNopiN2T7xw/wjAwrfdX3
1qvluPB5cZY5Dz4dIGWyey2flNJk8lnVKRryzwSdWHPRb3m7IUFac9EYTJcLCr+VImP3yyXFDtIz
dIvFHpFJt1WGhtfEpYjxbOV99XeGjVcHZE5kqTL7d0oqj79d2LRGokc9gS7mdEEaMUIFrBR75jh6
htQG6RjPnKPrxI2ogaKCk8wRNmjEahjWRHHnIqWrT4o1LeJxZKtgj9NJVK2d6JdLGG4dCe38zcC9
KTfl4WOIAjZ/nkRVCY4Men1d1J3iO7CLNauMhm4M0ZEBxmAu+GvDgnWtGQ5v/8ApM5XXkfk/9p4d
8Y4KSCFMPoPnwIUyCKqKYtOpxthPqrAsk2K3UKkWAuXNXSMpAtkfXGwtEyZ8xg/vakInjmhcmx5q
Ho5PLtiQI8kqpidlu9KYWdhl5vZQHZhkJ+W06LXTUhwClEfctlfYKBj5gq/8GJ5sLtWBcrsHKrGx
EsXuferVJb34eMxEQ3+eVV0PuKvc2NjwOQbMkrdyMlZ5uOeDQyQfd15RbcN2VQ68lpgBTL3Apomr
A7M9Z1ZC9+UNNzyZCMKIyEbfJGMI8ShZEOpBQCe8DY7RGrjBsYWSj6I+KvGFA8cjwlN1TRjAwGKr
fT3oKll3Ez55nQZGIpZPC5Mw3lALPlHOpQ9GyVgkS8l8egi6c191KfZiSx8IHtfhKqJJbmWUPxvU
oLJC2Da3sEnSJ5Ssw4nDMfsLBsZ8wGg7k7FaSTqhR/dUdAj4I2R4PZDxdPTgzzvjCEKkQ+4fv2vk
leUqUJ4l1BZ30nldBIHlfWqp+kAexWJMUN2/igRFwshvwoHalCBqxM+uDW9zilMc8HZfhfm5dnRi
QPSLGrsT+Iz50IAPTtKRqum2sLx4DO74JHXxwI6SloDqHIZbttPkarHdsMRRrSj04TRRDxco9OU4
Muo1bgKTfR13pjJh5SWUKybaiUtSV+vkGG5DefOS/EMHP0vqYTknOlo0ojIlcg7+VYSb8xiKSX/p
+qDG2Z3M8OQLnXN4/zrW9va5Qpu7QaJPMZcudhHcu2beYeoHD1Vj8UhnXidCKI13HQCsHxp6VvmK
YkuhSvn9AZwbw2A4TlprTfm3SXVpfAaly3qLzHWufaoXs0VrfUddxuyLl5WwjnnEhfWVVrGQByCq
uNeZTX6TGuwGCj8KOM2WAjzIJM0Vs8bGBooYzNH7yFHTwjxUpL2xXKIQlJ6T9R4GBUrcOEGdo15N
k/CvCdfGEzh+EW79EknlMBAOS+/tGC5kQP4SmSq9ZoP3C0G5Yw4uPU2MQB66ayi+h6Mag05/17O2
SYA3hak7AiNzhv8s1ugIITjOHx/TCfXjxcGnftGM7wMfDs4qeBjVbRzMxVzXEYsh0Fw5Siupxkwu
VQuqKvbz8bZq14I0KHgbtR4TLHj0ZgXz2/pS1KL/YBx4ow4XgU81dVE6a/OfO+O27Mk3wwLV49GN
Hou86NYlY2jYhPF8cEqtASs72dkSyZGLR3Do5/6DbLxJzhWkTVY28I4UC4ajH/sq+xCCUyVf7Lq6
INtJUYckvV2nsFhNUGb8Eo/2uvNUEQBzfoaiYrK38/bp+k0JMuab4Hreyo3Ps56zkh+cf/4V0IUl
+U3D4IuvjPcLWrpSo89coXHVU/HxG8ErDNeqjcJsxdME0e66eA6deu6NeWw4W5y7D4jCFsycVKV5
bcW56Poz4XxVIZQp5bGOzsJu72Zh56oF4FugSH0ZaTd/CaTrASvjpWuzZR/2E1B9JCledq7gyTTw
4U/5ykID4CXVck7PCldWw37vyyjR9AYOdkm04R73T822M4h0xKvgS5hl+ZXeGTxoH0cuHE1H/VoO
cqNWV+ziyevnjKtxbGwUvclpJLewGsPyF3hotuQ4817hAWEJTAkOsHqT2H9HFzJGQTNvJPITVOZH
PAMcONz8TgSV+7iNBj+NN6dgIlZQucYTH4jQrmqLqcBydPPrJOev8SpSCzApx9FJG6Rs8bKjno46
HxEoCFfBh/yff/ECPwcTmt9AQcXT9BHBPft08cG9QCb0HN9K+A7EDdApbZTn9TnDYvi+iZ+turWq
X6Xc+VNzZA6Z8EG26Xnu92H5v9uskvSuNc1flFBW7U7y5UJX9nQZSo2CfHRfxmv3ImO89Jh5okKn
6eFznM+T+KBOQsTeLdvj6LlnPDrSn2p1eYIal2dmaSiJaclZLkBi77chs3jTNYkHStavDM4B0q6x
QW/JH4xAwhwmqOiJGh0Beptc8kx886iKeONaTasD2gX7PamSfy93w9SkCEsMe3X70D0r8wHG7oGf
eggjRP31HK+VU6SB1vDKtPNDIOsfk5lsQ3aQtzPrENleI89/CL3ZFDQRiU74ZaEUqfExIplkK0Yq
1e76Ul3Y3wtpnnVqyDnWGCBmJ+/TDho8Wbqs/EdQs5S77H+wJaxgOMimxXPy4nnmIX+wwBvHpwN8
G9OZ8q6l+x3SXAND9INJR6O4bKWMxnt5KlbpXZP+FMFFiwk0BOb3vgmDxiS3P8F5aUS+WTGn1Rwn
YVElbSKB0TqDTsC+KB5vo3I38EJWS8CnVa4J7UxS2JEEPcXSwpzsTlKKKooVhbOKWh1H3FHdHLE9
Z82xulLkWZ2wMT+MtY8vpS3CTktf/uetT54eAgiDCI37FIyR3sgZnuzH7gvQomECi9rKn74pVrPW
XOINQZDNU8pMfGDcJCKtQNF4Ro759cYaWcCezRmX4RQUs8sMYpjk1X8Qfv2mXxrcOutBHJGNpkXr
oNMvAEJLxMvXCui2uhXXiZtAYUIMvLfs9HXB2oV65fydOtmEzNpBLKU1KrxTFZpy1Ow4Shu4NMcE
iWkPyCeG+0FPQGHvJO57Leg9p3pNI0A61YcSJmIQttEVZX7ZjaUookcMQcLVAXoUq780ti+dxtj4
8sB1qtJf9vsIbe2/58sQf18rIWF6NgRslnTVk43aMHlsSGXvLIolhiBs2Fypnkj/ljsZJvNbTZ53
TJ9E4DyJAEFiKskBo3A4SEKc744lnCN0gieoNvKcWQ1vIfDFVs0IlVGYZmGNw3yvt1EWlrBOAxDX
jdORNRaDpPd4imwnq3nODOp7So6aRLpttjg+RwQI1UwnrtLLv++lR+Mn/2Eua31qCCU77FL3UE/3
NQYAsFX+YhhJd0F3aXxSL7FR2jrC1HD1vRXKZvWBU0KM8SQvc01xgbiSeG3NQgNv58WoSEa2y16j
D84UpAiOYtiKYsB9yVo2ICS4jCJdu3XlI3UwTMXBpY5+aTbMyF5P0O34uJB8rUzAk3Bhz9JGvf4C
BXTmLx9flWq1Um8uya37yD2EDOt0h2mqBoSL2zWKtcB3xjdR53zWVAI4ye3WLq+OMrhxxbvffDQs
FOCs8AsCbtHWs/Q0DAkH/9K9BAZbjvyKt2AXe+Q5sBaLp6kS9o7rAojccbF2kM2fCS7HNqr45UKy
aOd0PER0zWjx2hMtHVFr76kD8jqYCsl9mrt0eVDACuA1gXjQN8wXpw7t2uwvJOltSgyx/nVta22j
MdWTacRKqhyaYQi2HFKnvu4LZBVQYGCULQcKGSi4addj7lQRKppA9t5XEatKf7RVnY+S0eddVzPi
Uv8yAPFMvtSGth9oupN+AsjtM/GJXbyu/8o/hhpo21tdIAyrOBBldb8PNlhvlQ44cXpRdDrfacgr
gVcl72IP6OLxUZGGhAzPjG8ggy7hJjCcxvA+f6wVKwVn/P4GFT/QA/xRqxDrSaJmoWdAQyHEFA98
5lYSgDUGebqs5yPq3kzqdazWcnMjqEJSlNst9/MlAtt1MJ6ITWKAY7n92WKWviqw0rrXuusrQyfy
JSYV9xjq0kn6BLUnCAlUBr0DxF1fLl4Dm8BrC++NQzzG05WCwVnXbkfAbYggZU48mSkFx3mI7F58
sffEWbYF662qunKE5693gGXDQXfiw9MNqLAIx7oBVGbp/UV2aSanf8OLeH6il9W70WYoTDlykdMJ
1b+Kc3bLJimUl3sjaUQYR0eg2OLRYXpGEcybzmg9DpMKIf7UFhRIfDb0bHvTrGe/Ez9wadxkgjSV
1kMc2TTKuSgwslc50St5KYFcrwAjrbdIyGOBvYcpdPMUL3Rjmo27Ra94QE0Oix/Cvq5xUVUKT7UF
uiRDUivc8p6J9bvwqmLYM34pDs757Kv0Zp3VTTscmLYXTmVNxcanlq8TZvT1iTUHcsxWaup4Hhm0
wBGg631EudTNM9EbDItbdIrygYKRBWtEOmJcz9mOG7trWVOxXt4XDtyAl0XuNB4J0/SPLEftxl4A
m533ulAkfyI+X4PGjfDKHXb+g+tOI0YlLsGmco8gHcLmTSGKnpcaVf8haYVgINBubLHsERFp6F1X
v0/UdeFszVhc65Tfo6UG8Xr/kcr2XScrTvytDmNKV+WfMf83m0qRoi7LT1JinqdnTkjWutIFH8r2
UZl1CrxkHJ/Wf61b8U1SxLRpc/ktCPQOH24WJwfS0a7JSrBIwWI7ZedBToTdw2NNnCFNiV1MOmyK
ZhIMx1PTYwApqv4ZEFF6sav1FXQABfAkaz6BrMixfYOsrVnuxSSPDBTPhCcjxOUB1IMGJCgyM8w0
x1vCnD9BqoDU/2Eps5JmKfVwJpiG5rLwmp4Rccua7fpRfR/hPuOCtyvA+5QvMqJvRpnpEKHFWuYC
uQ1wo3kAhQSrZEea0FEqjv6P8BwTazPMXatYa2VHieuih9Ut0YooESnHs5BCgYDUY6KgolJMwsxD
eck0PmFSQBKnmJHmaGNRlIF+SiLzsRwzKdR/yiPOOl1+5V2QrYjMlERLJXptWr3Tuygek6fwENSr
gdxPnzXdDC2+2p6wzACRk/kp+6Ef4kTSrw2mzxtI/sGXOtdZiGeWNBaFJwvzMyRgjW/QJ/2dshPp
FXd9hwswi9i8bBsfZBaW34uLd9Ho5zvvNK6LpULbStFJRCu122A7tkirCybrex4+JDzH4a/6fxt6
ZKvmNg2hfX4dMu2bARaZ7Ra4ZyOrfDn6wElAvXdR6hEixFLScn71N/OW+YAWDkegeTVqaXyo7rwG
3j9hqI52MMnO+uqOhMWnJjZeMFtpeh0drLVj5v1EqR89CR/r8rf6vFrMP5GFqGzP7D8sT5YrNhn2
u5vxBPJX0ihN13lA4HCsthpZ53QY9bCyveNAlgm4sIeZ38PMFGOQ+uxDNZeJmyIODKMJmpBOOzun
XknDga5Ks2PnzdIk8LeYarxrueIxOj4CyKEjW1sEGQYQNAmTe+mHYiqhn6Ux66kbp3O43L4uA/tm
NX45jSRoSMHzXc91TGwHZrQrvILdFqAj7O8asK+a5Ai2oZEX3T/z5rExcamNVf8ZXIBCp8LJKqQw
06vODDn/vcidWBngfJk7WDUkPzfbBYnO5zqAAfjpQWZmlkFW+xTKDklF0ZntWqDQE3++djPlbJf2
hurIDIJGZr9XCM2aBHsByTQ8pMIqzTAlgvlus150t6tZNQrGhbXzHoJTrCJIM+fGoazpH76OWmYK
NrAahzL7l3shHA1IYeh97gMrV/QEDh5lMj0ZVNKeMM3tzgZs1QEUt/IRxgjqL7E6uonE229ia0wH
b0z+nEZEnI6iuXdepOi2/urBH9FXfDQ8MUYTMumVOgutEUXP2PtuwbSJh2vUH1FUHHd3CR/87o1q
g2cGJNgrkUGEHzIO63U1yB9cFhYbsb/aIRGho0N/SIlf6uj9DYTZVBEnJmu7B35Lpr9oE1yc13Wf
a3w86tal81bUB/VuLZSauuRcNEV4s4yU8QqVJwkjvLYTtv7/t80TIX+/Ark/zIrzUZI4UakgQo3g
FqqjTAhDQPevCE5WLiRA5VuY0fWx7lo82dNkvU8L9pURE8l6tGhuW/orA3YbuGaLdp9uyyAbkQkY
rlik/RB+FpfRj4pMGgiccagzHsUZ6rhEw4sq4PwKYOhsByN+pivPembMq88lhJ0fdvSjGjfaOKb8
7mw6DKSw48yiFj5LkQofxv0yvoGUqNWM+BLjhmjwgBFtnd+qp6itZntyW6oRFacSfi754sN029oy
EIAMuGKJl8usSXgiUJStbq3w9VFk1QUgGZKs4z1VoPehGviWPcZNmffVCvOtm9PnlW3mQ9gzue5c
xRd3QKVWoZIkMPCLtWbPn1rgU8eeGsAnlViNYCdPBlSYAvXrDbx9b3ji9B+UK3tBOeu0vPkElE3D
cHNqMuu+yytCChJWqomZXqAtr4T0n2K/BwVMSbKFj7ql5b56tuAQ9eIlS3rqO3Dboe0FYO25vCbF
x2X31F0hd6cQ8WJNWT5PILZjqFeY2gNGlD5OMKnO+q/MJ2pm8zloGou0YbpmmQe7fSN8IKaovgpl
YndsGr9R58jWUJptAjM/yyH1E1Wyb6URomTRxFt1vkfCbf9exJo26nb2YlaMBah8SPxRzmyYXi4Z
yCtipC92XXriWxoei0tEA1yKMR2xIA065lMFmtIiJNr9Mnb6jenKTdbmzlKipKybA9ZoR3ohCJRB
/+mEYalT6xP1PBs9tl78tOUogGy2k4Lz2z/gJNDHbhyQK1hwkVuBr6qR3iJ7fOyX23aGUoDU6YcX
rC/rsOAbk+muhKSuikeZ8Z9DwF83wk0raCZcpCwPh0gaZz//fgvw2Ie2CwHOwsWiCYyWh4sTJi6f
OQIbdxYpa1u5CIKMpea+tq8+EmWNoOX4FM005om0B7SGlCbh670kF8mGzOrKHVm9sQ/ZUb7fYsKB
32E7cjFbvlXhtYhhyHv/46PeUEAO2QWa0cwNVTnFhcxx9d02D3G4pfnJX30VxCKJm8b4spqVFruI
mcgxUQ2TZz8X4aHorN8MqehRUdTgJWn4NyXCBOv3Gnr/1Q3wPwkOWVEd7chaHaxyoQA4I23tt9n3
T0V5Yph8hRpN+NBpanDmboxLV0g5oXHGUYjfXRA8AuMXMxvx752JyWXUVag2XhwMimFuZeD8sLEV
TjvVqmxkgv8qEEEdQlNlm96CT9N0wX1/9GgqM7b9Atsqnqj8zAaY+IMhdMCDFsz3ulRfics17LwW
F1DzrBqfGOUDC2SZxZ5zIrLiSrAmjOJIt/bOMT3C3uDliEawXLyQ5CqRjzHBlCURK4EpK/6vLBLz
UXQHkr8K8HyytjMM/u0r7+bYa6BpA7YiuUbOY4W4Gi8onR9wtqjXz4ElKFRjFNQJlml4xh4zOuvl
u1JJ+1k2LT/7aYaAeSvRG5tCKhw91e1Hl/Wiz9oHmZBAPQve4YSfcbPQIHlqFs7pYSyXK82wAMsK
TTmmYqzkc731+OKvzbciTmpL3VTw1/GmqQ/jjK+jgBj7Ut3MJyqSrZVaLurECou+x8o45fCR0JUH
KoM2G+aVlhfc6iU26CdCAxLhedab+LdYqCADhSJX1dr+tEDS9ss3z9/kSvdgIs1sWIFwld8hepto
U8rd3TBtkZxlbKS9BEBflDCEiFwR8N2tI4PmWBIhcwyKY8G60FHQ9xjhKX31YsvuEakwMVDqkDQu
QxdyBttRkfoCt9h67CIskkSK9vAUZWRHlFKNiU8tdSpr7sybENM7RZBGJrjkGmK8Afwnuv5eiWVp
HPf2h8x3dur52KOtUohFO0rPUoo+hOpUe5hhv29Hpo2/x6gWyRVKHcukl+UKN+kZdZqMJ+qvtRpi
RXfGX+jlguX5JH3imGTC4BfILHxzfBjP26E1ZtfhXLmATmAapZqwSu/kRw0+w0W7lQU0JitHklwY
4ef8Z9+qwhi2nE9mEjSbcaXwNU69k4ig1IIGFNpGODYJ+A1xeGM0HK2RT1JkSb85zVYVZzn4PUG4
eRsXaBOeaYgQH9NwEJ7oZ8hstpmO3pNgI6un330G1D36foUHWLknNemBjTHYo134vTO3ZIHYJ5Cn
yIXVJ1iFyN92YSgh8RpRogHm2WwrYPFFN24Z1yQyBKMF+1pAL21Vk5sFGWyl6FHfZCTCD7YXp7zc
m+4/bFSUXsAd8fqyzyxbBgHb7yyD3PfzvFjzQ+ddKbXMrElD9+Rwj5Cj9ExFNoL3ScRXa9qHrWYa
caiKAnxuia77L+NXcaVldBdcR/wARqkWkH5kmZl0mvBO2lz0XzhL/eKfk9mHNzEFOCOM8Z5Rvawq
VnqYChGffxJ2VZdN7yORGdCrRfQrJq2C4KQVMrqcpObX7VB43VAY6sc1xRCDCPMEytJoQ/9GF8aq
Ro57Z+Y0bobb0kJvW8CDqXjd4i/Z6md6UlpCSx07/hs1WucQ2Z2Sk88vicL1J8Z+UpnBpTQr0MwF
iuwfW/UxlUenWfHxSKHz4tgxneLDzv3ouNCc9TSWH2oo5s8wX7rxnqVBoE5vKjmCYYPgjVYuvObV
24H9Cg4fTin6tC8NB/ZCKVUg10lnaJl4GpeH1ZyshOVo5PlYZtKMlVJ5v6QFPGYk3HVWOQOIPrWv
+b1ictMZvgETvmHt20FCsvFDH9BYZC0TG9NPittmmXTauG/JJigNCC9ttoJ1eKcY3IgQkaU77GC9
uStxB6EalKVPP8MGEMKjVm1WQwjLiCtr/QWIWdfYZXpq84wOAi1cZoO/dGXdkJhFQneC1s2A08jN
JSZGNEhnziW7BARhru4mUyi0FUhC1GRHsLa7l5yxwvo5l0LxWGfpquCE4WO7E8LCBzjSRjcWL44Y
PQW87zCpgMpOGyjEoGUB6JiGOEfxdxHajF+8WT6WLzUb02oX3OHjoyvbdsZP2UWTmwbNCYj4vWoi
/OHiOxgVPnyVwledYK1uhIDdAwNWxUIi0rvFAIGwAiTN0u1hrIHC/BHRwJcxxFYjx0sNynWdZhIk
dBLYcmmIRnxXFicQMIG5iiUvqLJEGyopQpmjUbGJ0puSPQZ3jxKxZIyXMFnUwnG8QSZ6k6wUqc3m
xWYx7foqoeW2jqTpW97Lc93dlec/mQynX9kTGfAZkKEBgGrgvfGtYAHbtLQCi79M7AehmpBUD4Lj
G47kyYAl5u2GWDxtebACmvxUPV/qRaPHr4uGBlLy7du4uOID0Ztxsup48VkW9P8yEkuGW3y1450d
m2xqFmlhn06hPCi62xOwfPd/IHsgQ/ByE89KoK5nvkgayYkuliRLhD3bwpC5L9Z/y0zcj7d4H6ug
kQDQnWy1AQFhD+wycBHgpzDsfk68h6TvydJPeItVDTqrQd8uVa+gWX/SQq389q6cktUWAcL0vNFn
iKzjO/87/6EEpbBgBPF/rJcvUqHvp3VpBulbZdqcMgu9ZdD/OpIiW6OdaBitkr3yRtmWHqj7Njj5
z5dLVYJ4NxlmkOLdocH/wtQ7X9syZVWDKzzGro2MrwggYjJGFliTzaVV/FvHLxsmUiQlyetB+mNg
zKG9gj8lQ/9u200qLEyyKnIJqYLtB/za3vq/Iydwp7KMhQir+DsyRgotBGq0M+/mG53SF+E/BfL4
GIhl9NXkeq7EjYAOvoVOmwyWFOcI7dz0Rnj0MlP91kVW59OZqwhfxRMSxbw6klp+1HsfHrsO2/1Z
P++kDnp5HytDQjkaXoGcurMYU/Qt69iYmSHQhu9+TJwJl8KiEjuQZHPFhEGdDlolTKAqHXqaaKDR
Zd/YoapZ2sC5oCescDtP2GQgYC+eZRPUj+Y0KjEuqRBLPpJSbWWUnuiVQ/PJYYkW1C/shW2ZwmE/
x1NaToGi5uRM9D1LecNgSQ6+QtJHPdPeHDSlAcILW3aCDVLKl5zj9Vaw28EtcdKj58c0ND/g+spM
5e1yw4GHNYrDbB+ObjwZANJlebW8RgiUrVYstLL/zI90DRso70dudUGhXIQR/tiZUcdJ7eEF5gAx
XdQvFwJEgsZU7ExLwT3iOR6rNvtMVJiD7wcCaSN12oUjpFnFSeqr1G9BkEJE3/IemWehVcIBe5O4
JkXefyw5EUGeEapYmefTo4V1SiO2f8zfh3M1zccSk1E3gBhaz++5Yx/xltAPbjuheezzSUNkXB7K
TauZwvsiluHBCkWE+ABE78GXyuAcY982nTYBBOnlpvjPvZBiqmfdbOXF20snEpMJ2ZxejnUvWAUS
AgKM1+8bHOWLMxkYg8FjzQpkkM4NnC0UH7C9eIaInjoss1MGhrlMcyFDrHK+PFanz5sVa61/9vti
6WdJ9cLPdGEAqtWicxwdIS5Y93t1dvwbdcqCDfi7jNTBYjab07N/2Oj3sC1/LJgr6e/pCGXQlxIU
V9ySChCXcUFx7l+XnHdycwK9tPuduDwQHavCuwGUBFAYNLBM4r4wRiBzE/si6sXjAmV8AJ96Qg2k
TXphCM58OTPQZnPqtIq17PBrzuxw85wtyJ4AehNeEsilNlC+O5ctoetv6q8L6pw/xi1HA44RFoRL
Ulz/96/HFcJRsVGXItmSs0CeWJnalzMmbIeZpPK5NL1TB5nHS+/HSxif/M9/71pR3xkn++oCluCP
sVFbw8/BLqwz/WJAaPAz0jA2AhZo0gRxZqAhSviYwF65hDoJDIWxkWcY1AzWI8R2uACF8xZPfSRK
sPVN2+CnskRAr3M8EASwVQa+FKk63DhdWtPhNSnlrLsUc0trILyNAm/K4rhmPGI/Z1odaDPjMurl
6ErkhMDfsQhpop7gD22bnhBxwyBoPXOw1+1dNWp4FTprWLtj3ik7u0Fy7lw23106c7XaiF15BV4S
ldE2JEhnMd+3TFWQcL9ioVFp51aNxCkamvqsvkJlKCtWb/MkyLazzgyTToug+Te/lkZnzpQcgHvZ
9e+dKIN+i95+XhaKtczkz8ANh7inCBpeC9zbWFeq7VyfnKDd3Qz1Yv/oBmql6LJOQY6ItX6CQMGt
r3JMkDE5/Lebxs1CkIUCxUR3QSYbMtoB2m175N/m8qLZ0hXCFC/6gxiykhIzAab2+epx95DAGTZn
4XO257mMFjiI0dRPn7kFYfM3aQ+8gUg6ehz62HOdb2p95OFW8ay8SBfIQv+tOheDv6Knq8OfKeOu
fjbpsriHCT91EBOg7LE0nGAkdR90WJGd8J6h88u+aj9xipk3vnHTWJz7KNBSiG7+FqmAZG8jAVQa
BAqRNwXr+gfOF4JkjaK5JKEq0CqhrwMlXBP2JPY+ATpmTZXmAdg9JUzElj3zXp5J0Rv6OgzXw8Xs
AF4DmaqaYJOMoph3h/kvWlQxAj1l7QIBIkAeQs7AzGI3RuetMgFdyMv0dEl7b10OoWm7boBGqHNj
RkATsAndxh7GmHqfS4BbAkml0khMFVEjReqFL+cw6u3ufteoF9c2MuoCP10dTQOafwJkKMYEyuvB
2V3ytZiNioTubgls25jYXT9plA4cWKrXX/C3cEUgBZbKXELieffwsOlWWeqzGMmtiqpRAotibY51
cYXiOq1w1sVmwkmbNhNbxvKwswaqZJI0V/cSZTCZ9KfF9Uj1NIjvbZC93kAol/oJZ8T9HQmB8Sq8
DtZqwefxDToP2Idwjq3x0okMS/50CimRLuydcknFrTyvnxaFkmRVVroe36TAb41CSWcsYjnT6Ujl
4Erqg264c1k49BdNSkpsrDUKpVvsJYJ920OPPkPZLnOIJT2J9LXXQ5e1K6w4oGx8XyAY0XgFVLSJ
QKnrVRcyyVGh4A1ixPdNlVTHfHjlH86OxwfUZ7CuQPFexs/Vpwv+eKoaezZ47w0I8bllv8J39OES
Cemxgm19iK9fwjAAjsh8FHNl14h0AC2cxI+xswD7ULTKJqI62A9HEvar7X8kUFqZv/NeYEntQWkh
rttVpOLvvAmBLbBoUaOPLzbZE4eZI4Ra4dSWC5w1iWXQKU8SKqtw4R0ig6rO+ngEAJ6XKAsnr+v8
tzZew2Le2xv2nusgBaJGWkrI/rAqzdANjnWIWYN1RtlVTXuNrrHP/KIw0l9f+dJg0uC1WLOeyibp
kfCCdVjG4sLq8+AKH4pu22b+CzuRTRXUcTGOzEb0SicHCaGB6nqxFOq3y//t14xnSJVRXrJ/g56Z
X7u4etZgFVReAStlHN38EpOs8snlWlvafnMcYSCJp2mIvgKamLyN+gloJYX3H0L/guvKEkXDcSfE
GexjIkXnvYjxPKzYlyT82A+cA6iTbcU5coYFBGkRBhYIi4rct6P9KWDV0NHZMOj7qLOOCTDij6Iw
8/w3FzgadyPg5yrO42BknpgWDRMiUV0K7sQGKlyP5MMz4oMaWXrG8UTjfSjkAI22oZ07o0zlfy3m
6RSzs/ml1fdhTqHm9e/dzkhEX7p+ifrAGhs5przzYZo172liP26sfz/TyEOw7WzrBDFww0tXPs/7
mjoy46h0gGGm8+04qPSaYQ+3ViJUS84yYPq7SmI5CcOl+XqamGc7hkQifeukTnvz8Nn0HRHREwvx
uloo7N5FO1Gjvk1LtAEshKt5U7uO03PUifkv1c6ipJkFHwE9+XrAHZexZqYOKB1hnnYS6d93E7Eh
3IeT4TH3atP/SrvXJocUWejWQbYsC+HK+chRZ0KcaZ9ibEKT49WPXmibIt5MRFIw+z/LYqQYlmPf
hOpSm8/sbBfeyT0LvDI7zPYkNCZZTg0EKG0whcEEdaIQw7ABol/VmJ/zO73WyEXk8lV+xlL29umg
EBIypLDmYh17grzXDQlDr5VIY2DdXyx/lo4B5NGheKlCWPGF3gMwnO94bswm9ZAGTyCHsSH47hRD
AiR38xfTyfqz4hqkwlo6jPRSn5GJ9MZBdJlriNMLAJVK+0iavFk/NH2kBQXjKdvH0sSsaF/Ex3OJ
plv4Cc5wExF8VYK0P+PFdFycoS6TUpLpC285Co+mg5FTQuB6WG6qXc2yRK/FIMvYuL6PGAvat+QT
BrQnkSrXhGKKtdwyB0I76h4mKmDqEiiJwr5sEjVioIIweY4hf/tjnup8pv9eZ94PO8tVoWqPzlll
etZznZalJ/XWsxaYqW5M5fnEQ21SrdBBeHC5JfL3H3pE9mmm3eYa77NZgKmNYKPPsU2a6CMVepnl
8SXML7OD9YCN9Ish5G7G9esLxGbxbtQe0/4Rf7eP8JabWBLPnRhmjZaY0QwWHMLdyknsQvszbbNg
sgncUpU+6ldxVlmMV173nNDM7EmrQn5sggi+hE/GxQnd85p2/zcUlHRbUbxDt/WRPb+kthbRxxoc
rJIzNM0sECBgTm1spKPxbiZj11vuRib4viYqaiAQqcgHso608lIq/lBr6OiLlioEHSD9bPULzUm7
y/uRMdRfdZvD2H9p2NNcgcPBE063+2I4DsEmpcabp8OtKOjQxDkkssnlE+ktWB00mP87n9rdDtTz
akCsBIXYNeuHN7MLszv1ZPGNJQ8lxKF4VG7rE8AqvCeXrO2NajRL5meWoxYgZE8kcVGCaBk5jkb7
Yr8Yuv/yqLLbVsDWzJ+vThutyvhcLZoFoLEB3Omk/akDa5EbqoRBf4iXL+Egs2HnMpa8+Qy7Jrc3
E/UInvpIMLzajF48Fn9bxJKHH8h0srFz8aTzXtoskilgzA2BjAvPyoY7FHlE4hYUsPX/CrBFVl+g
4VtKKBRFsyUeRbgUGiJD3d9LKx9YVSwMIkzK8p9rZne3p8dUA7FUVynlhGeBLr1p6tuOW5EK5IrV
ZSDxWIxLQrR8vq1N+uNl2wq57j2DsE/4uWqZ+GRsjOPb5xqa6pifK+EJ1jxda971ONFMi7qUwUop
iQSNrABHwi025494G6d5MHkVJn5bbO8c2A9KPmrDTImRI2bQf8bfyXR588Anmc2Iz6nIve6LgFZk
2r5BdToTjHqaS4SYclwYehEW1DSBDH+zK3fOoW8e+Y5VrxUIl9U9HQ0pdLqNXls9wlylBtEdITNr
FSz9IwE7ba1bGmoy4N6kXcUt+FUNZ5xGZz1ggyC8MR7gkfj+2w5Vptq5cgwbhENuRVx4zsPJGN/c
MEJtUglM9YLefndkAckD8aNLwcUU0EEvyjPpIlFJlXmLb3kWMQKcNd+ZvRJZr94rJpx7IEfiVG0T
u59dA5Jrg8ATWzSriWbA+ILyvXLAlOtqD4bFt39f54mgVOtRVMnN5Hsn9Oil0HbyUZ26elMXFUwt
c/lRdEo1HVbF6f7fCHslvT8t0VXYusihsl2hGkEiMgeRHxF+otYH70815s8ZG64tBvuH2zKhx9WL
ieDjEaAFI5eJJ0nnMGJNxpH0AGHQRgdBHSvLw/0BjNm/fKEqb4qJp6l98bVXC4hmd9lwtLsYnKsj
cv68wuIO/yPJbcEiPerTVv6pmAVB1rqFddDqbyNCOnQOf9MD7iDjEqgUUkL0eeZWh3GvlaSohnnW
hf4+tl79lH5Q76TjaFkkN8VgdgIhjztgIhDBrDEMo4LV9PUcc8y/xZ0XF5ztfuH9oNctvkGu9BvR
P6cYrOFa8K+TMod1AO4VGuHzoTb8csf58x5iZciWf0nEHYc2T307QoE1MqVJPstuWllVTa6jMgAR
Ms5O8mbIwEijtqY3FpTVPTdvnBJFmly/cqpC/jOyO5IzJWJvTUC7V710Roru4ZelA0LxmOiOb0Ln
C1WjCCp3GkcpuWiJjwWjw7HTVu5oi42L5AaxR/jkjwYo4hule8Cm99PR3lh8NPGwQYA2kL37Nx/y
YRMAfC2e97VMWnpOcS7AmxnnB6kaRb2OVnGDi7mfe9PUThev30ds0TfSY3WUBw8ZH4pgYmZ7ueJG
jmwVhcNAia8uPIO5tdmT72/3XiosDcUxADEbmUaNTz3YTPxyfFAji8CYXXp3kigUWmc+Jly/NC2R
KWog/hMJKYdv2nekjKu//4skrNwht+8tBMIDF0Lgmr11mVL+Pci9Ve1tqNxYhqT0zCRN+kcvItGz
EKAKtByT0vc+htBIP+acmhrKltYuvpCDIHk/+cMUh2KElKUe4CqsVKchVzRNu8L0nVcbjKsHocMx
a5CDF6ee4tYJ1t//pLbbIJPeWPf0SXWVQGi9Zf2jwZvpZGJuRTPwiOFDeLD84v20HYPKY0Utze2N
Va2X2yVOoKGN1l0WhAwzz5ymsZQKgBbBSKzdm1N54nxuhjuCL20klg6d0sRdgDBAU//FNzWbjK5b
zwlXXDx1i8RiebP9l55Ep1FRDq7mzkBeDueY9YAg2pinA2rdiSz6vlinmNJHoaIiwNNUaTHnLx/X
UaCJOBCDzbi1nPth/HwRdTd/jLIeY/eA+9USBjw7JL9xOWjlyw0rk8iCP8emS7r9/Ada1OBENq3R
5Iq7ERZKypzIoytsBRx6+IdajEffjVzE9jBR7D/4wOz2saoPSJ71nOWseqOIEHzILtnbWycu6EdQ
EP2FPX+F8j3kueeAlQvZyA+maGuaZSuaycxehi2yxeS6usvVhpoRvWkCbMZji3PeCEWDpwkr39kp
YLwfXbeCZRdZqDaNj6VqPVCV/Nfpwez5Wjl8JDjHNppyeyCCc+69r8FAOGm5X8MY9CLhChmMnsfu
Kd12dN9mbLKQZWsecNFyZZ0RRA8w6bcs4YLhjoHR/K6vvAZ3sV/ZrNJFGENcwJZs/utkm6ObRZ7B
XMMaEj8s7z2K+BQ/P4fv4o7yiqxO2y+z4rSvLVbbAf3Lz1fmWhFY6pfR2TvkvZkyyqV7wjo4FTJ3
3K+Ly0k+b+rzGw92DlhoTaFcIRyvh2LGHTB5JE8DtZGbVzwPe8hn/3sqdHLohElvqj429jbhaqlF
xCM/EkRRjoJ3nIbnT5iUgltgFCvb2M4XjlX1lN0KEqdpZLIYaFlORE/M0cDzwYeV2V9hrlJvbXBV
c5MsoJeEGmkpfg14jkM9PAtQft+cUovgcOnlENioFR37egb+L9sEYyA47X2APQHubaOS2E4TYPtJ
n8ynfwmkYtGnm9zuubBWYvKceVaj13KW56Lds8ZTS/o0tMtI6bjC8IfxUhBqAnJETz2SJv1veujq
j3ZShHKNdnfZ1jhMAChpLHHTiFi2AA7i8tsRDLLYsSCcFL4ekn+ErcyC2CpqQI6ZyVpWyzeqBbKK
y7Z2z5X8rqtfhgamEA6K8zew8q9Vp2u1+NnzzuOgrwGSQ9wfs8AhTTZwoE/FowD8OdQaOy8qfkMV
87OBZCyIg36OZQXlkZxi2wXGIqoRzz99lVINsg9gKwTQcJ7DzINMaWuDV56YP5zvFrblsnXb1anY
W0Qmxit7RHJNvGUxdAj9ZHhFU046NhcuUBw59FyiSsbHWFwqdLPXStq1vSYbnnzKlUIBTyhoFf16
Bn+chiWtJJZp00S/+hJKzUk0XhI6EN4QoAB+9ut5SR4UKB1b8lhZ3N5bj5NcLTu52KwEO1h5nyBI
sOvX4lEQIGIQXGymxr7GDidAuY5da5wauV+8JAs9+liU15XYoAfcQ0UM1CPs4xHvw8h9xaL0YMK+
OBqbAQCCEO/PF7MYC5qMouWHoxFTXOwMrChL7W+ZuGefmnKU/nBIjtlUp2dt36iOFdiy4nL3/3sZ
0OrFpRumkUVgE52n+QPlhGTkl5DaI6qZzm4lLSxjl3FWIr+19CqFR8kvE7M4rtOUihLROVXfgcpg
GhiPDTSI1NC7KVe11I1p/5/5oaGwlIc4Ze4dg8/DkkEcfb8SpWBVKLyUXu/IaWrXul/cuQWCo3dV
mlvpjTXNeWpVB+P1W7qCSqqAXKKSoyArSJ/yWcSzrg9QVIYgsc1NqnQvkRIYZAJXEpf+xsMVdrAf
Ce+Zh1S+k3qUJ8d56tfAzYhGoL9PJEfSxYVHd6AP0Q1KmViVES/GGu3iH0OAa8LDjoJtvBfyehMT
qq5uEAqrNSiQ2VTCWnStJxsDsILhBSrcMsbFOj/NdHgCUI9dUAxUGQluXG4FIrXKfliK8fIdJ3ik
Xi/bNpmWFzJ9ihv2YGgKhJkCIfJ1uXDOUp9nN25b1qHCj7bsLaUDws0xjm0JmFfB/GZu6TK0X3H3
OX/guIgKmt4biLjw2hBf2Bt+9iMI+dLG+aC9+0pEFsnLBgdN9VDjGJLriD+ImIE1pXF/t2d+fcIb
6MH8ibaA9X7sdzfmJZl2qkkuNMj6N2LvZandXbmV/HZ2QsbZhEMMaTsiWdmZax3LZCRuctuFoXe8
Dgh2B1osC+25EdbUlVAmPc73JshuSlBi/1qPHyB65CS9JBIacrUQl3TNARTrc0QeACc0eD2NxS4p
DB630rhIJB0+gq4vzaaBiyY02KzRcxVoU/feJ53kxfFhu6vHhhY1HjDg5C3GeF6VtQiaOdVQo2Qq
l4o6GqYE1asswglaY5IYj2mkkDyoohOEGLEvWhEym8o3kgr3/kaTLbZcLUAGDAuDX6YPfinrZKsz
8HHMQU3E2MP850Cr8ggLZ1MFwKRuY0io+hCP9KNtFtOi8FhTPDh202IhVnpzkhWRLC0cnPkYaRIE
1HHRl9HZYsL4eiffOZXz8l2Uic4+OS1tj8P7c6BfAxZA3eZ7xwpVwNRm6blWniRd2fFsMTVRumMT
T0EwjwlHxOSOGgl9KjkmlRgBhjcrA9Nbc12ePaIao9/yu6JqgVMgtq/wHYdb8RYtSHbUk1KlZTL6
bwMlScw5gGlvFZ02b27q2H6lkpT2kRQy4frT5xivOjrSRJZsi5UZeEpdN3d1Y9ie1I2PPPw2fsFV
w/a7jAk1Fdj7FPi6H8aaC4/i/pZoWNOOsRUjQMc11me3GomEj0qtNslYnS/nysZVACu5pvmwCzpJ
h4HVkeDedjfa1lr+lH/rado2qDZ8DX4g44Bd+yOHlLvAQiBbGUqBzAPGx3BaDZkbVs3E0qt3fdqO
ieRxXEukcyQIMxAz0NOFKPUlFLWcalVqhNmDasG2BPWVyBRpSnMvKT78Hjinme0Gz0jwS47YQp4X
QXgmVZrLVTOUL3Rc5yMrlXMOF7YcoKubTlJic7MISzTx1s5qSKX6KxHq5TqLNnOtYT4tSAkDWXpz
Eod/ZrgvgZySzk2zYZyAkAoh/F/QF19coxaDyJM91+SSP8yCbJs4Ps2h8b9pE3ghDxp5fYSquDg0
wpg86+niF2eiL+0PLubZhcRCLicR7WeJpNNKRKJ0iIyTdYIzP9E0lfKyuNypb6Zfyr/BdW3R64Cx
oXDhb5TVhRe5IyVHBXj8qipDla8j6TwS+tu83tfaiMbwfnAjRWzEdNJHISAd4JFRhhAWE3JX3pQM
5AlzadyppnNe3ZsXc7kWpYPyPYepsBHUBmq+um38FUj+LRQ6M0I0MIngxHWkWG1pop9O8R9xbeWp
DaTkF4ZMWZg8xmjdL1Uw8xsrFn8n9iMO8Zo6lWSCRHXf1usfYCd3KIQJY6sIV4/FqNqDIY4kCa1g
pogtJt/1NleZdtGRQEdwnH8xAMSl4X/6eU6IdlI5EiNWAKNWR761li1BO0Bl4MRRtDAdubMfIJsp
BEchbWKRk0yLvBwTsAtESsFejx/IpeTVXU6MZqA7XAi/5EApMXE5c9GWUDK6PWTcgKiQx9QmgJv2
rZOj5KfLc0sSqzRxXzL3xqxZ3Mb5Vng8hjrTqFO7eGQns0QGvLYk6066/1e1rBrM4VUvM8Cu/LWp
HDCaIGFppeZ1Q7WTKGRqyU/1+zDOKLAtGzvbxeHDJ/SPiZsT2rScw26NEfLzrXUm/1Btg8PWZNOu
/zzug60u0STRsEKuKlnXm/E34Cl6JFuwCQSmTTPY62Ir8Rrmt7hoUuBp9iw5f6ONcHwj8k8pKs/Z
StsdGrLF870lxRk4nT5HyUeL0XzKW2axmNQoEaKrD1on/kHgfBDMOIDnUS50S8ABuRq+Ht/JYzRe
1tGA0oz/ufAiB5LsrPJ1IOwjesAe27i5KP8ThxzW2ZsRzUBsMDNUi8eIcd3/h5CWoTiGoaX0/w3q
8rV0uyxO10ju2Nw3SjoPx6B6gl9HX3R9rbu8psoSbmC7Je9SMSl5FPSc+ptmOmB7Rvr953DUxjuF
KOaDPd24UDbI0ptcMfV6idzayDMIu+82oqIbQWSd5avem8pdMKoPNIjDcrw4rgKOeTNMPPrZWxgT
IXl9ogqOUJlFyAPSSOaonqn+fDfn1T8nFr7oo4IbZPSzHbrdqFYvQEzmTpfwMVJ9o3RpKnpPuTsu
kJJ9xSUrF+XxMLZj+8FI2ZWXf78bK1LxCSYKXjyIYCJXfcHLNRmIicPUh9PunxqDBzjRrv9Ugdb1
yg6xEFD0OLhnEk4wDg2TaU8t/Ar5SzNvDNkb7eA1wse6TwLNArVIEYjLLXHU299GjhSf4rth/B0I
PWuPxHoOgFMFAAFaF6d/y33Qdq42UHEy4c09jef7G+o6d+5WTzRQJk1IEPJpCerxVBkAdtF1Tcib
xa3pXH9BRa9Mm/lGioM7n+8nUR3fbldUzdQs87kb9C/YR0eQXSIgwjNeRQUdXvQzcFxu0dCIY2J6
s+vxhMPWHvkJwO5bhOOBlQPOq+UCcRSk34mdB5ZiqhRabEcVtcsDzJNdkW0Zr/NaEs1Tebdjxbvo
mqRW4MUyvcqP4+pzU+FyHyraszkV21Ay621Mp39us67O+EID/HjN22W43gBZbQ5BFGFZyALzY0gN
Oy9evDpH1hrgsXsaqPh0fo8vbnkrEW3iFtctovPu2kDcKKSM2C3DYCp5zu4+vl/hC+6P4uknJTzY
2Liay6NVXerDThPmOgmWTw8Z50GOEUPmV3qYNOl/sDlZ4Ewtu09imL4BoTsIMeVx34I29zOx6Wxc
GE7OWPC7OFwB3JxqvleQ4G+vBBUtStQ84Tzn9Ah16bYF86jjDHGu5r7GlcvA7qRjeJsvLvdl1AOE
/GaZTFVEoMXHoGqp4ZHWq+jq/JHj/Od7kECknzEjCHBRF1Dxoe+Tyo+1jgz0R81dMVACZZyjFVt/
AFQdvo75giZWw1/H2YjPqirIVcrC+5gIKBJyk81Dj3DyCctwT5DVkphntB5NBspzi3AIW2Kv3kZn
wTxu6l/TDMHoCe6xwem6H1cxMht/stAX+YBPhYB83ht8/4fgS6O6AqRoMhozbSPXNaQiYEvlQUhN
FUSL2eY2itsUv3n7bFNpDl0PDiphdgwhOlATG/W9l0XcDND8ZJuy9Hc7SwbI5kRkxSWWmfJIH+YS
UUQH9CRDpJR9tei7mLZpbPXPIOYWlJT4W2jFL0QJ91vhdfWzibPUn5KQg2M9zhbYd58K43hr7VaL
ZrWwJ6HZFgAg9Y5wADwWJPcFFVvO4A0A0hY/qF4rQPunmYD2ZnCev8ehejQdG5tN64IH0ftwEpfc
Tzr62A9Ni18d6I4x0B3FSK1NE7YJ848rtyzuUm7jxIAQBfutNicbw7MVkq1XKkozuuua+4EeM1en
BqePzoRWoberrRu5qmHrjN9ctBa2HgjbI5csy/tr2KQFNd3QnZTDAzh45ZA3VA8XSoOEDvYQlNqd
Z+Q45nAbgaSVilSGjfqBrPsHgfsvvnNXNWPTDmCfU0EZXDPyPaPIM2si9kaBS53avPnnDrJ4usJ1
OJo6wgWKxMjMyOO6ZsjKz7XVoVihPgHbhnVV2DDKyJnUT3QaH1rcFmY84RLFOBeglbS1/ddr33VW
f0/FE1ps2reS5JvoqjAHTj/eeaDA4azjLeFMExtQf1QBXBSTpdfcMSbHOdniNKPEPOUf0s5fWtvO
FFYDEJDXLKxD0mLI6HEj/v65q/wVzACaAlNIl33sgoHpmCNg6NCyMjDsUFxKWV0LYHzWGMAZtZxo
rNT8xU85kIVSbElV4TSJfZGMB6x1lywf4lqGzyx7uFtcVAd8mvJFKAyOiXrpwB+azkPiUKgOSsST
qX/KWsPjQBZH5OVVNeaTjlKy1L+CL+ABm5tpVEoiPwi2b/Z5/KKdk2s8sDk3z87AS9U0SeP4uej+
2WzqJkkpRkc7lg6JBK2OWkOXUqb+Fx2zaG54TvBVich2IH5Zkt2GfNF+Smty5fa4znjASAb9ygRm
gamjgq4nwCyL84gZYl51PwQicjQIkbbqA/T5SK8yJyACzDebrSO/YLhCNOz912oovu+ovA89cFtG
xerveogMHaV0gU6m7jjnAwVjEU0SGdHjYdywhBGpxkuTx5aYM+HbzXvaccHFLDltBtmqRRrFGALH
9ZLHtEqYS+XeZSwh9+gb3HQwcsd+LsM9fP5KfyuAhhAfTNZIlSwWZaebPCqVG9zAz3i9cZ4lGiHM
ISDdVOnP8SrTAW/N+J6e5uF7yN7OqLFse2RGLFQ/TerQ5lqKyVw7kPSV0obUmFLwptNAzmTWHMRi
VMiy5JM8kzoe4sOC5ASwNKiB2KJlwkcbH1sOn2EOsAXdYEy0SivFEK9bkIAmUut6oLLDrSYPTkCh
Far6QoC0QayHz5tzNpHmu7Q8tSx55h6oRW5RY5457KuvfBbq/vdnbnGXtJPgTuNiHCbLkKI+tfDW
A7PK8EaOg/Qd+U8+0W/k3JGt3OlIWcvt9JkmBTzRcUFLyLQ2x41OYlXvvChIH/TCmewW5lCJYJtL
CDo1yzp6duKoLYpE9h7px4Fb05XTOv1gHEJ1/Jy6KF0ogJg/2cOyxadN3MTquAIXuUYJI6SulTZr
nKQN6qhoHq1ENuEbIr0DzrGwVrf3dPnDv14aYJx/3mwzDMPuIE8uIpu2f7dLCygGAaMkmUzFUk6O
U4oIe05+0M84t8kH87SJLygiSas6rIQvIZBfC7fBsmZVayg3FH8pj/tcnZo6KNHlAPPhCUQ0sbNk
mhU87dcgzBQ4BfaVDM0lxaKF0p9sBtjiB+pPKpHpdj7PAd8+QQgDumogFLbRuf//S0whQOZMwgac
1JUjuvH/iFWojy1T9kfXnsR3UPSUyxbtNvctHgfs6lyoZ3aJdJsMVNaaRojTfZfwFBjzTidFgbFt
+dHkBqa2hyp9bmFX6gaaGMDH4M7Wd+CiZkBRB3F9RIOy2cUf5ec+6Fv8YRG3hzQ0aP900k+G9uoh
UR2alg9QzhX9LSUv3i6+5qwvgAkIoRWTlnRdp38DEI1rFNXpsHZqrEy2wYuN+ukNywVLMD6ZgY3N
g9jPMbfc0Ejbnh2llAG8JTB/6iwmEKjzmE3ivQnzenBovRKSM0QiobmIjfvmKPtOybDpE+IL8Aey
gaNYlVeHfv6FHhisI6w0ME6zlYdYyBk0UQG4bW+evalbfU4wxsmsOZ122rC1e5DWpcpTIMZO3I/e
ZgZQUUnJBrkBUjlC5w6YzFuIsFnt+shXtGK/5D2s1s/ZfEHK78ZTESbJOgXU/k0kKKcm3Upobcw8
t6/mevkniHK0Ychl3mjCsS2bZp6w6OGvpIwDpFdLvo2qNcETG3AW7kTTYvUQncpPeZO7zTjLf9Aw
brRo5FNjFok3nH0T5HPop5kQ091EzQX/apAmOgtZlBh1yxiTFyoDiULvn9GvswdoIeHu1Vw8EAVt
i5Ys+RI7wuKHcmOderdnD6lYlZ9CKwzboK371pz/UkDb83ClaTjmUeBcy+yZD4Xp8t3tLQGVQ9EM
CeKi8zNAsEcL0sMR0pB2xwcFVoCmXvQYZ7YTe62VEg9AUqcZwmNdjomvfioSSwGmvXJy84tGchCB
u+4wjuO48YXojcEFfLJMdKCrS96pT/1al9rWCcejnKx8r7c7jvgQUyjPNijqnR1GiDLFe8QqRV+B
QVTAU9EnKkCsAZt6O+B3Yl+mF0cw0wgZxRFL7JuDk2y7JSJNp+El2h6zrKjq7kCk+1toucMXM9PJ
ekyPf6Yi2asSTnVQqw3bMvGWD1tISxhR2KNqKC81gmPk54VR088IWnqc2nRTzT4wv4qDNemV5sWa
MwY8i1K7+HHcRQjg3NkZ5fhGW+1NFr9y++FPl+twzM/wlurNHiJnz7OKLETHkQRRbrQ+6olZICRY
fkPWu0FfbzjaNTFDjPSwTyrybuhQV43rjAKdZgcMaStRcsqAmi2qpyrPuO7mwE/JisB2b9KFP9Pr
RPco6kOJaHM4sdPktsYBRNsTjL3etN5ZIouIXtlApBzgUXCBNE3/XZavPuxuc1JK6eSQUCEq4Ldr
fOJarEIa1xYuqRFZis/9VdnH5pagfAr57pVVGtFmrhQuePP8MHL5DtoGV/h1LT+iz6G/mkoMKZlI
NGkmeFDmHDNfrntBGG7x5+6K1VwI5LpNAZ4WG+lTmW7zAi74CEtr6uZvP1AQVD/dC5YnLDutyNEj
uCt+Ink7NeazlaKL2hBNPvrRdBfixAfQMzeAVVaTS8PEfoo9Ey3x1OPaqrke38gZSHjxVXA3bQeE
4u+rMD9ZBY45g5nTz1sd5Gx1+SvVpWIqLgxAInaE1U7CQO/Mxh4ldEChv9V2M+ZTxE5FHqTabq0z
FEhDfT17Ha87TirszcN/Cu6KPHmg5WvAVaHH/cFnAgplp+yhk/SNdm9qIR3B64NxiJ0Xwx61J0bg
Xq/khOOuoilqdCPXQfke7zZoks/CIZbNSIJR5u0qcPDQDYsfSMJuvgvSH4OLVzApO2TtM3EjX22/
O9ub4sS7CUyCqjYEdbTLAXG+iwRhY5cAiwqR3vBvToejDg38y+A8i2iR88E0IffcnOSHyYIpDu0x
xXg6uS4xcxPxKzqptcXOBg6/hbFvWUruCHaIBPrZfxm9sh6/43mrOYtUh22LYEfZLa8tDDWP7Y1a
UMN9mM/0AWmG7+aC4jxYizB7KoSdJNeXzZ+nqKQL4V/VDfCPqBpg5o1ElJeirdlGgi7IqoK5/sHk
VNgcoIiaFiCL+sw08StZYI5NDDuVuMLjJBShnmOJymymuL1wqPVLq7U6qTW51X2MhUTd7uZ/f5Cl
BHqh+h9vwhgvhHe0Z6LyeHkmWjBVprAsfpyHosInxavOlC45P7mfNcd6NtMzPYeGTmEoFaoa24c6
KJaNg788xYRuttgRowbDyAQPnYO95lPRj6er2QKIPHU4UzvlcE7AJvk3tYOwt+Dx3r9ecQNYoIaa
BnGK4p+ulPl8KL4o5ltYb4p3r3sJISMWZnAHLk07m27Gcx1WXe9R/If4Fxp6vYEbcQXPRKvkA9aN
2n7pAtauPO6BZ4xOLUjHLTsIDsa2CYtvWewY1oXQiDbbdXWExujHMK4IyR62GO+K9S3i4IuU89LC
te9Me47lOfhsQIlqv2EWBxAD0RU0P9/3gnGZxfyIjRQeysZN/WgnR+yPSwc1zRrE1J6hiWitvSWU
x9/h4GIwcMH3nmBMzSI4yuhjz6l4aIP0QF579Id7JuOJTsfQuILK3KroH5E20FU1SS7aa0mnwxx9
IPT8LnPtd/PafjJp6VGSF0kEc7GcNUAimGHX2REQXsxewDQqpt2YJ+GiwS9aQO2nXST47rsdyOxl
iI3y6EeI+fE9IDddkpIGM+9UmmXMuwi3ybIuELJYxexbNwcVC2jFHrfBjzd87jbVRqCXORYjSR3Y
yM0eCgXqr4libgLUtmRHHGPtJui9hezV0CJZ7EL++FWRNB4bCHyo4bXmhYQSOpTQOy1dITbIAteQ
27zp+4+WfssJlI0UelHSrn5T4OatIxp8YCegClW37VmL+9X4gcyrLPdnJcFQsvlI/UFLnbgkNU+u
vLUBeYk6NZZfvrrNlPp3A43ZmBbDoxwpyb0FA3WmiCUs4Mnh/JtZNlLxLEuptYs9FgiB3MlJKGtE
TG/7Onw7bN5a7QEFXD3NngtyOv7RJsPCEWWq2AMNK4lB23mgg+cT3JSPxfArU6wzXDGTQy+/7sMh
wlGNxE4QYlZEwsqKYRP1Vo3/wVXcaCf7A8f4oYKmum6VKxEWhjbEcgQWAuDCsnJFnSRaGbPCIVwU
Z+996PRJwhdOi5g2UVo/Aw8HvnA0oMfTSHqgMe8HY1cCxUCJYgAt+uUvEIaZBaw+gIiCdijs/Er2
HyNbb6c+Nx0NCJivQAiaMgppzRiCXjdGncQTOzdVhRFuTfju8+PaBjCdhBDfbyyKTBGan0+ZAeLT
Ip6frTYSACPMRobTh2+91ZuleT9dfedMmZunCVZBEGyZJnLUQh5J8Q+KAEY4dSRatXs5SJpR7Wuh
5D+Nravf8ilypey+TqimxtbHkm828f/aqgWzDhqf/ImnA8/UKqoDThpPnDDRdeMKBhcqjasHkPbu
AEbBhybuPSYX7gYvqFUEDIF/wtgYeAYynOi5q9K2CBNpkZdFekUO07b48+/qHlpD/sc2KwehrJnr
1p93Z61mQNO+Yogzd+EdcTXExoVDJTtXqxPeJzGporGqDJLrfjQP/xBgRYaadww62XbnCC5n8JYi
iiHa2DUkEz4ii+DJ9mYaP01tAhsOmb+SPFSixLZA9h7auUebCfdrRaub6zsqkYmW9dk82VGAiVtJ
E9yaZaaAcxNvZepzcIST63M5S3jeaittdvBaErSVMFsj99x+OovpABvHKjRLHIaU5NBphne1juxl
3IIkJ1p3hId4XQNuqAEhkOIKALZvElOH6S19PCVH6qAqUAGWMbwUq3xDLPsYs0phgO1D9ZmbKAd1
bAGrR9SHzvfhv/pfgIV/FJwa+JYt9T+77wJfaRavzTROZYSYfqVmWcQSmCL0P5Lpn6hetPpEro7O
np9jOglPpEGXk2A3JmdDgTlQSLIWtVXVBeCcb0hczG6cHZNp3HsVoJN0xJ5/e7PzkOFOzp2Eb4RN
YjrY7fqI6TSiNl94Nn+s46fqsVG+fOhUt4fJVkSB64qYds6iUNk7uCRe2TrfbsvtI0TEwgK7UlZf
P6/kymD/TKRqN8gYOvwUX+xmH2HG3pbgfgtOudXSRMgeoNBI2nzwsXK+4sH9pIlmieLCL6HnbLup
BbxTpLFkQjoHM3GnexmRTu7Pe/rivhBeq4FM92sPQNQu2qV/pi+HT+IFmLN7W+0Osxd1NavH1/M3
DNdYMD6CFzETvSrOIs9sBR9ggu/dg6CrNR21kdLXAmf00z9AuYeHRPqwiF70LuwviLRwak0VXBp7
DdVLfHLgkPbgI4Eg8GN0K7/wse1XK2B/u6E/7zf7BZLSEsZI3y4XhJ0PPuRWaayAMz1qsdysT5lR
Yuri2UMZpDExj2BYX5Qe4K7qVD3QMDxNH62aYrt3+DplkeanrlBPvoehxLCOOGiwQLu7mApsgFhM
bX+4iFryUXt2rv4VpdJSvKUesl7W0MeX35QYqlA1IBb0OWypePXyUsFEeyMGVvBKctVYpZXIJVx4
/TO3wFqsiYVqES1glDzFbyyLszNNVYANyCuy8JYy5tQWJSJkR4kIw/yok9oV3T2u200DDQdqAyXz
+4LhWIa2orlk5IcP1aQss76hbPWkia9L19JVv73X8O6K2YfirAPe7qFGYRE/KjZNovXw0t+vatMD
gMKJlMw6xMgGU4jjhL48P3bFHWvLf6chBUcd003MrDe5xadTvLmCDFyviG9ip8DXF7lb+Yi6sABx
9WDt4o4kXXiARyXxIkzNyUg39H+OfU3DYNVn9aSAGGkSAHOElBjfeAxYuomRWRwgTBuWVag94Li7
jbkCu6OSGbmOP1Zse4lm67aLBVTon2eb1W2LtCWsR8AyMsb+/YQjGtPM7ThEk84gYIqpcdRsTPJG
OgQqX7/LiCAL3LjSKo8qhTdtvrKogYvQJdwpr2RqpSS6arJWQ90+96dAA6jt3pHxlseVUiz+pMIV
IGrqAVwFrgZ7VCcUSZsD4etfMdn/3NDWf1D58O5Ys6yKJzihDYVgsWoHaADwLo3IlHUBK4GAzls4
vUdLsg0GD61v/7ocyhrhSUZ+Irra/dj8tuaaksMOgQa0iHG+74vKmLdqkc/zEplWgu2vLCkEqyk3
UB8fuDy1CV9+0Hslk+zuKiLFwmrzo9PpNKDkoogoWmC72Nbz5T+UE8LkhtkY/VjMQmxEpvh4g2md
mSE/7xGYcGKBmdndQhED+rvUllCwe9EPS6tioRDidi/nwu1N6JVjsAxFoLivj6EZOCEclpC0Nssv
bc0zvORSsYnUUGDnkmsTBmOa7bP+JNsaSuEzP2mlrnqYQsTYftrtn+qLg4A57cczRPbflYSPLSRT
+KrbN7MoOT2FHchgLp043Vk0V7AptSN475C9MUNa8vDqdZ1YngLAj+VErIuedSUly85xa1GNbpWj
Sk/Y29Zk26tLW/rc6NnvYe3bufiUs0KkwDL0a79w1kwqRvvaYTwHWvp1w3euUG5SWdVifs0huebk
JaPeCQn+yHVYZ4Bzgjdki8QLBC9YJ5ApvONe9J77wJoRVW1lAka9votDMJUZ1f0OEam7g1mRM2hF
nLPNvlqElNUSqo8OxwEqQ01+4iErvJ+5BeaaFTO+JUDJs2fK5k3sZn+q6pM8Vna+13lDqMx9sWqg
cv8LQbkjKT2aCH2hTRcAl8Ea9fC5HbvpvDi+ZHNFjnfEphoq+Ec7IaUK4LmNomfHPEa0NYE/d0+n
NbslkuHqzjf7JI0K8fVXB3se+1AxNTtEqcMPvE6mvmfGSj5Z0nHFamWtSKiajkL4zYKCn3b1didk
DuHyYbWAHAfud2ZawDpyELg0MrYhDXCoX7xSH8mSWlftNcqUKPcWM+IoDKLMrktsNYXmJKRWua/H
Y+nMEzvXp0SrgYtt/7w6j6FvJp/9x38MkOgNBPD5vPsuqwbAk5+ty49oNHvWILyaZ7oKVmRQ/X+m
s2LRirxZpcwDOzVLpXzlx1F6ENOiwzG5yVmt5jrhOVZqY/e5spMa4d1ifTvoW12vm1XK+ow0F7W1
V1jUnaZL+cjqnC/qSIP3BZ0Z/AZYb+Esb8aXjMtpl9ZR5bel1805BW0+Q32VwmipObV/l0XZW3nN
qQvbv0eByJJ9TjfuBDmHlIz7S/9ZugV1abVJpybTnr9I0P1KWnnG2IH/XX8OABMRQRsMyZvN4cXN
qYxcWeA/6deuUCM2gvK68CLV+Wq+mPu2imi7Uf1uSOI9k4K3nMoEVwYEY6F1Mht5ZSYl+5CcMGef
TmWdT2WTCpQSuVM1TGCYM/xPqgaD/mckVN0pWkysRn6xY1epK6Z0GNi8HiJLI+O01PF+q0DcMzy9
SB477ChSbrPfs3/0R+XFZ/lY7ZkcloKEMFHGsSQWp1bS9iWxMgHYB+xE9a5F8ObxkZEwPqYPgtwB
f0zbrO/mcWfTzLdubpXvszzKtZNyfKE+OHIwTS7Pc2hPUUAu1Yw+5i4eEhnoh86TG/OJgS2vVJOo
aexp1jKbc47sQQXycqWMj6vVUUd3oQknhBmzIiRIEzO73fQhavUcZwRbIhbhaoLzaC7i/bSWV+el
db5zWwBMeBqzaW+pp24bLrZIF8j/3D9Q7jpnGXOKXhmGk957LtZDciR2mlrvf9qShNWcxPzTMPdW
1qrWUDMOiM5tDRiE87e4Hw8fg4PrHQrwtcs0ux67RqyOGotkeiWfzOkbcT0oqbxdrIY91fUe7A1L
xeHPEbP/VmSKHmA+jUahzBAecdC52Ph5M2pUtqqqd29NTnlkBAh5+ZiJnvLRBg5TMu4E+9kJj2mi
AHj6nEQRdFbnrdHLt/YXS6Kwajj+Es3kAjlfWw+CbtzMqg7xY1AnuJtO0MkEQOaFTCEunsMfbgv+
5STYJs88Ewa+7nRrvct1ajqYlNxqpeht4pzaHPdRuh2DP3vh0MPth8DlrjI03Ccz7MPvydAPP3fK
VBBzAajxKPxAQkxAp5l/2Gg0MnoZWOTOhV5smISgBvOlSG3WLAPIzyxRka/aFNXHTHOo4S5YMRw6
xtFSpi44I/i+3jPNrEPeelFiJ5dog2cs8pK737+3rjiU+x5UV0+YuKE42VPa874MVAiLqqcwly2G
5YQ26OmbRIGIq1Y8e08Jl5xOYRGNBgxPjfMRKIXnMjOVbSqI7KF/n8k/LbOHnRxTFjxLvi+/E253
iVKGWOL+Q7JYwan7X8TC6R2nO0GVXuwhcEVIZ9wmq90b6YBsIBvfBXclkUUWGnkrRrrwN3bu2epr
YEj7IAT9Vam5G+/b7IE6ULV8hP08fTAdG5tcB/IxB1WotM6qPGJS+n9DqnNlIRdm4zvW+GzvK5Rt
8/CnZ6d3wZjg+ArTCHXevrvmrgVP4moHuFIxlYyTxmOOHcSz45MJxJr4v+6Ff2UmGSB5aCe5QNsl
r8ptlxvRnU5uBlQEYfC0Uxr+bNJ+ZG0QmXhsuTy9FPcjpQJ2hkTXOs+WCenJj/v2X3gDylyw0jPX
/O864m7WSQr6NDVFKNjzDDDh4RLaa+6qflMsMp8nqqD+HhVDmAo3M2a+lRNJg5hYnuK7hFLb4BKB
QvEu7weKsjw98kYNiY953LJ0TW/0BBkbzJu1Xy49cb/cHqVm6Y2b0utFsQvv77bqp+8DL5KPcdsG
aGMRzXcQ7McEK4Um5NKeBNeEEfvqWy6NUyhsAF0/gzZppqi9hEPPqz2aOcEE3yKG7lA9iH+vPe2E
Eo+yzZ2G4yN4blRhT/wxHKCUfFjpp0mysoLmf1sVVoORDQaE52uzJ+uwR4M6qnaeiq9uyHA61U4f
GpkCyIJGmtyxaRv9CwMw79X03McsZUxLt4wLTLAxOeYsbE88zSumhHSxPQSZ0tK9aVhnPGWYd7Iz
ZP2JI6L11Ba6kXQaJH0FjIr43rZ7dqLMP0wC4gDMvJzoHrqbmXRyD8fsVOKXZyRHs1PpdjvmGQjg
ADT6uPZ66J+F1+Ufb33KL77LhxL2juTBfK3M+CDXmU4BImJLCi8LnYsqa+/rPu6npwPpQ5XOf5kl
g5zj6SmSUJI6kp18scQ9bSk4yOgIeXLxnQyxf+IuuaJ0qRL5rJE4MwCd2Z7O/NmF7E9jrzkhHjix
UTobxF+YhiUuCj+nuDbB00RejiZRdCeRxjSYxxggZa2XUvvxLviBw8c3THm6UYE6W2pLK04BbRpU
khxWvEkPkIWOcU9lyy2Ji/mL/I7FWb6MWFOQNnpAfdAtEWohzy2UAFiwVGXurIWS4BdTNDidxX5S
1vYy0/WP35Uf54XnTFgCw1Iy06Y/68U0QS9SRRF98LHo0LkiFBR5f9SKrY2RzADdgGR19KlF9ITG
frdU+kjFLLuC7ritHOFx6cf3Dn0QNXw+QF8azUGrBwMP9L9bE9VKwMi7q+o83dpAV1Hyw75oQI0e
P94KKMp2isSMEpLC/S8JY1EdRU5AQ6V/CWTiO62xZmIfGPZa2hjHlCmvkFwJ8FYajFVT6WnZUii1
8czWKaAq4qWmfg3f+uJ9PbAShFrBqYMfdmef7lKAsYjkxGY/OJnkFPiCVOCGmj1EcAUb7OuN95/d
KpSKeVUEUnCHycw3eJ4aVio9gumNaeP7UJuH6kTUgpvl3A7p1ihVPgRpErAjykiIrEdEHaHD7eI6
EZKf7+ew8LDe9CmdbzNfaeBlH9m5c0wuugObxcuIrHRXtcWaT361FxGa5oTn0UUHNhHZIjRXZwvF
d6dNSlx3eGm8IT7xs2suh2bmC7bK1vM7S0PUzyY25rrBWbOjF82OmrYGBDjxOSU8Jp8EzDGiy/FJ
Qvt0y6hTQW4NKMMa41B91WRqy6fKHjaHKmqmOMtaFlUIR0G35ISqkLWHVR5/rTEWwtnn2e6Z7O3I
xBu1Vi85p2YH9rqLPE9CM4P81n1FNVDSJ1kiveHvKsoSg1CA9x6/BB03me994e32mLOOc67LVfab
DOixwplFUZw99of9Nw60YW/hfbBw7ElDkW5L0A07cg7T3nwcDKGzBeGtN6U9ELjhSHrTFISVxoPC
H3R0J8qCFOOQzMoknkuoh4Yotn1P2Iik2dvZfRdTBbSTaY0bw3ss8c9yv7LoYCCKaoRzLXF1rsLP
CQ6806ntlZ43trI0xQzVeK10QsYqOnTG0WI5PoOzX33wnEcY5PZZB3EDvNSptES2oppgsN19daZR
WRmm1uorT91g8rE9UmBp8FysIW6t2KchdSM9k5tj01nGbmT1wA5y1mp+XozKURmAVmMagGMRi06Z
0IovezM0urUCjEcrC4KUUR7z76lYMcswu4L00O5C6yRWKdrr/AdVUweFFaoU0ZFrZSvoYK+RD8f4
q2NSsB8bUGED8vnO+y3lUyU/CdRSAo2uYXkpCne+qxP8vFRI9BBY9w/39b7tGKaifzCy+ErQ8KhB
g6szJOG4Kfg6No2i6e1cqj6yrTKRiSe9Znc09D2SdqIIf3HjIXDC5NhFUIa9W5kxmkLOTriRP0Ek
+JGcjtmrX/cGElXgEFTOf5mUnZ43/JVVYjQ1cePcmWMxRF93oc16STIvB5+I+khLxkFHrbTD9EYU
gpr/04OvV5ivovsJw5EOymhsFrYOWuAMQ+PGnToSSmTOxkMQM5mNwsDMClMKb2XmLe0QhmrmIA2b
7Kpq21aRCowXFuFdPj1bugr1rNv9g1GeLAwFTm6HgPyR0QfTtcSjWFPmzNtBLynRAdNu9+gxnOX+
gg+EE1zXaxV4I0BGTjy8YZqG7fASzjUcuvGy+jp3HV2LwS1Fl0eMDJJQOfHDDW6CkH0hBJGMw9Wd
65UZnKFgjjtnH0U49wxjWCKBujL52S5BAT4mZJxV8PdzhRNd0Gpt2kl/JDwSA1oSUDtvTVMKPI6G
IRXxEWm3PBhW2dXQoQNHjDox2KjS23dEYufCunL3Ww9EpDo69kKKni79LvN8BiASRp24PS+qe5PL
/nre9C2clSGkedjLCaoK18CKnkD7M/p1fhMeI0rtzJjoyyTyQbYAvXEz9vrW1ea16jGGlACfzmSy
pkWwVq2+sRRNHx1VQaR7nLeaDa/u0YaH7yucLsIyzQiazqfCad8YBSwwIZP3mFQCxBIG64hd2Ndb
OHZZutGDvbh4wq/g76q7wv1IVFNEM2uKF9Sa3zhz7pawQf/DeNwaC2rgJRCU2edaxknNAhF2W2Gp
UckhA0ZfSTcWjAiyCRmgRdWGhhmJe7MKKiUd+1+/FInpsKD+z7v2pV7ey9ZEDbWqBhzc70M99PN9
gIM3iShGuxPSgvuxIh7wD+EiDpfjkMWj1v//SlCkzHAZTiHlI5sDXseqbjkeZ53UxCM4JLKBF5Cf
Ywxyalnk/pL7amYXP2yroFq78JCTipg+exIUDL6JaCIQalKRotPPpJ8w1BrIeyiFRmjPaVsBviZP
UtK8qmaFc+jjznaUt0A4qOqB9270mvce/3UDju+2X7srP9zodatgV/jfN6oPlEeGCRUI78hS7EG6
JyjqtzYOYmiY2BpiyXoRv+Ooe0MzSXoXosowKgkOLbMfpUIQdyYQm+JBiq6lfVbatMnmtlzs9Env
t60+cKvsC9XCc0iANBbI310KEurLxVLGiUI/R7o0Snl40ZxRFFm6V36DlX/NBBMfrMRR1Ho3rZeV
OcSy/kqmSJO5uCscIOnmw4bOC/9fl/N0Ez4yWEAxOyYS0UvsaRjjbJipxX79RLD24UVqEnl98RXK
p3h6Mb93pAq2ZyLmASWLzrE0/sZ9CxX5HvYBSJobF9jNd00FcPOizdBW+mgGfHfOWOLGZ5CuKywI
t4Qk9yveS0hjLld2LXdONGFccludAf5+J66w970aMV/DaTV93td0XB9HY0PkbmElh+m7djKzNQDt
N8Et7RWQShvPv7lr9vKM2/WswH0msVBZbzs+R//YpaIYvVge8eeW/ZYN/62hWDCm054MjGRTX2ur
OLLnbC2RmNxohfetzLGtXNl5m1YTOV9wGj2MqgcvvQ4DrpaHBFdSUgIcVNaCl/iC4ydNkBXtpujY
+H0z2MgDsyuQKPrcjF3YrEwtWFWOuJoUx6qTvrb9gQv5plfAly4JFMAHL0D6mp2wxebwX7QAibG9
VChMc73nC1t18iiBnTFrczlRIAuXvtLA4VEjxYfbmVU7EQNyYYuiDpXfAK7bt7dnkzD5OXpiPp4f
QjhRR9Jsws8l9EgLo/e6jpszesonUmi1k1Bxq+dCPW6pLSSYI0/eA9RXaRQMOvdBbZHa5CINNbAz
b2CUelcpdokRet/gP638v1WNjOPhi7uNKuhavd8xn0nsnff1wQfkt0bzkP0o/J8DW5Yf/Q7Q8ewd
+CSMT/Yc0Pi1ZuWI0pVGe3y+C0mhhrs71Jaso8boeaAkYcV2kL6NVRh2Mrn5SbfCm5NoSg5qIrki
oAkSl6KOQgIvOuabOFVKHZxNiIQlgL+s+bZgEJ/YAMrNNtED1npz9i2hRjyM0EHuPVP0YL/T6DiT
NsItqt5dOsCJ/cdbhKE2oRRpOhzV/B7flZ9i/sP19riWSFbx4BDVyDusivLVEZcFr5noQtV0Z8lo
LtX7uZBGyVzJ9e3VZlKur9spdsnKIzfHIgftujGS7+Vx3gVPb/UIMsXxfjfW0oLz3MwCeBODq18w
GTNCvJONkTcrJKTwf6HSs7hG7PdY7Y7yuJyow1qRhex62m6bfKDtBbSaTW04GL1eqe8XVqKB2eex
4b9ioyR1RhRbJAdbaVBk87UTHsujdE+vwVMWVW+aX3Pi3xI2z1tegPIj8lFUaOLXI5+/NIN3O0Dq
vMB9y495CM1NrbCaHPBDyq9vZzrS7n9W7ayV7fKh/ThXNjJt3ikqBCx8b2HY5Yejs8m9ZqH/URIY
Hg+wLQx8M3IswjM/8QC5Ln2qdA3Qk2LmIG6rJOrvf1jRjTotwDPIO57/rMlQfW60EtlMMhFeCP/7
pKjz+6zZXnMmwXqD2yWX2PsIsqokNqm1wJLDCExyn43J+7GbxE7x2TPch7DOVmyLVbt4P9SpFyrJ
eRDX7XyVGB5oLrhOhMGEumWOZTp4ucym0Pfh0k5yIoiGvNURoI2qCu1Ork6CTT57wV9nGP7nQuKg
cwVeOMAQ6T4TxWjCrAT800+0glYHkwEaVrjmIrE/SCm2MrvIB38522da18a58FRFGhngtFgbSnBu
UY9VbAgVriB83Krk7N3uBjei4NRk82oD2ah69lq/JYE2P6gdWNZIvJ/bOhK5iCzbX7A203HrhOaJ
H6A/svKx02h1gULbp+uxj5XJ5vFo7Tw50t31nR0HbSlRrMhDXJIO4ZHZ580Ju/ZAC5Wzc0evPTSD
Yf0vS00gnHRleSbnKenbwgTS5TBSXmW7bByxttQDFxZdNZU5W29hFrm6V71EAJwMLrmeTkqGxVks
W9KDo0fTaFnoe90Q9DDi9h0M3tkz1AXg3Nr1sU5mIWmE+C2ZYfTD5hY35QcYn3/O5CzeaR6Wyicu
pgiMK/ubX2S0wfdCx+sW3HYmoe9pMuEX6vxpVnzKrPQUSoI6vU6573IOZq12/R7qOjsMFWIJeoru
3BkVpolxO4ftKmTNXJAyHHKOA/Y6Prx8Lm/bd19RNzbtHxzqUYV87TBMw5Ma+6Tq900JdgCMKkel
9vpm9cD6m6icTQstezxL5bJjDHn+19E9hHRTIp/aK4PgdTNDJRcB3fMcCbho9O+o6PHOlid9wvzX
LLw7MceMgeULT+tswXybWns8VEe4Xk2MIGQFhVGorxb7cIkeD26yYqhn5zHGDFDJux7VOnm9moel
Kuqe9G58/TcsK9a37/G+R3oXl+iT/5HOvyGlpzzAz2Kczk1kNKJYT1byIP8w7woFiEnHPemWQh+/
Na6Br2HL4hEAbK22QFzOylvJromLzBiTKira7Rf6RJYxa2QWC2SxXqkgPDanpiCNcSoEOIaWC1Xd
QxdiLokvyXkCGY+iFjwu+/VresnV+zxGsx9i2gHpyGk5kVkgjHWCBK7w4WVGo/EgcGkzu+wpTWz/
aAkwfrqMAcEoIT14pUoSVVcmMmVPMF8n+ikZnGeaxEIRBmCYx84bNCseBHuXRvv8ZjDKIZAZMQXs
KDxR1DHDxrKjAKXmFjasKQh2K2b9qBOThiXgwl6A4P/P3SttBQXH975UJDDXxyvgAGIoOI9zvh38
Py4jT6AEFJV8Brban4+fy6Ubuj7sxUD6dmNZzsIQCSrJwMzB+IuJDVqTSK6AGf/6FH4ZRG+s/kmg
AqLICdAUbaJ8uEKtAIu4sCZxKiSxQD2ES4euOTErmnwF9UOD41mFAp1b6bljTwmfIZMDKE9foT8y
WqZsNknxGup1rVH+tHcUwtWZEySJjKK6ACI1DHyxsRwlc53cjsaIy1dvOXwhHLUhQIm4Ke04nqZH
JqnZ6P9oc+9dVr9VMoJH34ChJgpnNSYkhUQRPoaCyURw2QedClIU2IDjEpfofHgmhw2WVcrgqb84
T3S2A+5Ugbaob7izNqYjzo8BiMJdTZRf/P76j9UdBDPp/CGvvTI976zu3y4pMebxeyzJwLyJyeGW
EOYYNv8sPp93GsYBgok/C5VMq83XhLs5d6Dz2qAeoKtTUlZTqnSPE6VVyS6JgK0jh/rfpaJ9sAv4
taU1vvnrOUKxMNmuyOq4DcY7RKD7dRIUqk/ZTk0s8jyz8b4HLcAVU7e899pNSHiOzHuR5prRn/yj
oEUXxWdfE+RZFzOAR32Eir5MR+arlZHZ6VvTkP4Q+DMoO9uAEDJD59mdhfrQ5MGQqfvkXt7KGvNm
gidBHtsocpXjVYnZ/q47EWUW9oEdSK/B+Z2Epi4ZyU2BdUHaF4ah7zGh1Aw9soAdJSK7K/Tw/62T
c6Xouqe3ZB+NA4MCEuiVZTK+Z6dRNGHbkMz9kGGR+GjGJZ9YJ8yjGxzQU5opeIfUYQqsjnX9YpaZ
euG9K3EC1lebad0NlHigINpC2tH5uvHvTiQ+c2/vqo2NZ857UFOKuYqFz00wZ6mMa0k6oN0hxL3Q
xrlnnNWJPkHWCo8d2EZwMyE2h1edIeLzZ9dV5SnMSURigYpb1iOIUFdaFj2jTtQhuYXwGs0x2SpZ
YIvrI2cTfL83d2RzkYdWOWOM9sFFPm0bxTJfIuw+yzJ42FEf3bz7HFfIHeqQSWEaOkokkW/u2hwq
FVG/JdHq0asIbMTDjA4CJbMC6rGkJzql9rh6hLfXp5RUNwpIBMaNLuqZG414/gkpcebAeFO+YJjS
3EFVz4lQJLsvobPPEcwV4uTzosrFpq0OLvmMZ29etntAFcd8b93vQmx7ilFnXBd+aAFnZlD0IVNn
76Kq1Jm2uuFu6ZRs5aB4czaKuCaPv2V/fB9Bb8naqqzKksVnDV6G65lHs4OhuxUVkIdI5Y363/iG
HHc+sSNerCvwcsJUKDkpXfAKHHzm9XfYuUbOkbNKTnBDvSI1usV1r8IFsq1ja8QNVHu4neri1FRN
vJRsTz3mb2YtD2nuleOEuqFxVv8+2RHG0XgCeGQFZBSxpWaOGZZFfZczgy1Ggjm1h/+ViHpuVlog
wHPR60+LsIqV8PpXiBTdOesvpeQWeTlzpwauDBqqDWKKZxSKVHYc6mb8aHU8IYLrAinQ8VOBnsnz
KdZwREYUqCBuXK7vtnwGwqqbSkmBZ+GUT8Amb5TlfXx37m1CV+uENFck63Pt+2LnRhxvHAELIJb1
UsdHCiP55W80K2Rf3DP+ot4OoDVwq4nw6UnuToAG7DVYEgrDVD3VN4FNCKnGjUj7R33TD9lQasYl
WhWjEWJeph6FfkKSm63SJ/8foudlZj1Q7XvPIvv78oeIrTNWF3Ox8nYxUV2wh1bymJ6Q7cnmXiCo
XcCMzz+IKWyicsU1ChX+myOPHfrAHftyB3SwuUzRhoLOjt8xS2jRjPxCllW7rUVWpzRpD+N2i7xp
KWkoH+bRhqRWQQcEFEzCiXQ+6w9odTh0z6W3uXv8eARCFCMLdZkKIMpqkVCZ3NYKAVPoWJR1IdFz
IG82YYHHQKhpQjNV5PdCto7T0C3Yz/SnYpkmUHGc9ZpobWHlJm+TemWuWnVC6Eb2XHVYZI1Nf0xY
5DtocgSoNH+kMzk+ewmhRUJ4DKDaDYj9f1wpHXsCF8Cw8OVO5/XXqElgpLOvEygNGfyzhUcqncZo
XfWbrpdnCf6I+L64jn0Ezg0hq+IOlilGsDFJb9kEZDTl9a4KTjq2o8J49YgHSfgDb3DC7//K9mbk
OUg/huj2lVCSQksbqPEhbruw0hAKCZZ1OSkKurQ8j5uTrXvfSISQ/lbu7+NRVKMdpWesXTJpnMFf
V9PyHjbiOCOoId5XWB/dcxC/LhJhxBGPSAIGrvl3S3fNkFhQV28XM8BYVGXE/sXTxuca/Ebr5Yge
NuPH3ILKOwXHe+5ti/+tKFHrOHnd+oSCgPE8jW0OdJjMShjI1w3ZtBtx07gjLPw/FAXW+93pbTP7
gjzpRHReUpDK0bi0+b0uDlrWb2pUKVjAQJpuiLY+DSHDCNtO2zqZUgzzoznnlOewa/eX8lQGFDv8
AtilxhvOPaOyB3pc9qKMrKP8egKOue6GVrOKQ/oGd6bfuIVWF3HHbZUTkDL/YgwD7jtcMY5OayeS
4E0ShREjhHI5AkdX1x1kJUjGBw6XP3iyg0Kq05GFvxcOzwEy3U/fZgowKJd1sCeKjEUxXfxIKFBi
EVQ1PEXmK/L5Iu2PyO2HE858o/C+58dEhzawPDqINtdH7buFh8PnPK0W4KRgGGpYPyhxyF8JZsU3
2uswYgg45yGXeHYM85L5hBpdIncVxM3P1wCzZtRYtvm2mO6Xj29va0aoy3y6f5oOX++MxnQEy8md
ww8kQ4rpdUtiGzkIL9Vbmn/aZkJo/DM2VWO9hhLv8Xq36Ede7JLQ+vhYcu6ppoWS3fYjJwXUKWYZ
xVsEDbnrnmyBQXmItzlQUE4gxjR8uei8ILCy/D6v34t4MlbobQL6VHatwLQAQ9YI3dGwfBIccA2+
NfPBMa5VqA1FzexmTAFn7Lx7r+n8v+Ld0kpQB5jJVbvlrvHhxsvBr8X+0uVWgoKFtHPtyNGNkYoS
SXTMEX/gSc38ogpL5NTHzm9GfVMqmTbuLEgCQ0M04vU1JnD5clSgUAOWfHe/+dsE3TEt2ukqGrdB
4fsdJVX4QmXBGekTw2yber+JqoNNtrur+ngLDmQozZzF2WAhFYCM65FYJeiUENhVDyRRU9kVHBkI
bTFaIfR65xtgluq2SvJsXQAWhrPRIhbuB7NdpeG0zSzHZ5Yw78OeIlEmfb4xrxi7hxGXPr7dYV2a
SYoy9G8iFHoFpaAq5TLwbCbi58EvR9KvtcvAts+RcMwWA1sRgFNHPJD6l4jjBzYWnbt6AXy53QNe
tn0PI4X722uhk5O2ewiDBJzGUipK5Hsgx/7JuJ11cGcPqo/8nU6cUpu9V0GIlQcIBAN6H6HyzuDO
NwNQ3pRYl5i9JPyugWUtz0oYjBzQLUBzVpAoSjOgZrwphz9ZbGf8rylursElKYAOQ4wBqE539r3u
JAzA85Qri20hHajX1tpYW+cxMb93P2x9dn1zp69CnZObAnJlHxDk7RO3NRWzm/bgB7EhhQfTl4lB
xzZvXv7KUGsINRHKwVstuaMShT6PhYfodbO9i6g57JZ6qGZBCVIVrzufmGz4h2hjNkeos9Xmp34E
8Gf0t8YVD4G+uVyYr6esdvAKIRXTpEtIUERRbTobsoNIIAmtblZpLKsTCuLCAS1+OVl/TRqAzR5t
iaf8ZC4IZe8o6yeHYHbUC/JNZ5NN68uw6kk1MniG80BxRgeuz9tjYAvR32CcL561Wg5lG7aKSmzB
4K1JveGjaAwBs66mlltD246vj1nXMlaYm+W1xPb5Ox3k4hlWlUc1OwoN/idTg9AeTDKkHiq23kii
A06BotpdYjZFIWpX86dSK4+wJZmQ2IHBf0hQaBTETh5350AD5VPU0ISE31UD5embhiPFkaB76lal
U+Y2Z41+hQyFmnSBzsB9MyMIwX/lPiE4V66tZnCz52tAGLfTFr6oWSZFzeGfe2Lfn1qJ5ujhfEb1
SFu0HPdMSiXo27YBQFuWyYNL543xmhBGP4urSbGTmbsrJVqRxLVJL9YpA/vTNjEwjmbi0T2wKvt2
36a+Jv8erAURHMdN1HESZl/g9O1kO7ythUwMnO+gqmi5sBkabxNCnMHYWD7ZevXE2eEWNX9nZi8t
9Ql2H2VVzXUOXimIUbVri2mqavezeVCA9VpHNlOQrgMs9Aw/1Il9LwSV2g6IkBtAyVtwcbtj2yp7
4rdlU4ZQJdDISA5O+uK9EONA479AW/KF9EFnw+kPElHW2j0VKMJTdcSvrfLy6ZZ9MGGsAzTlKCJ6
01Rt7hluQ28gstrPg2PqG6CmN9hUBqwzX0pJDkrh2dy179xJo6Jr9OXVcRiDS7IYAbxlcQQBNRNC
PD63/ktMaL9+UMt257aWD1uyN9eSbK3c+Ht/Sn9FRGDEFqjH97hrfx6MIVKnSJUa8zjwLFGL0nCi
2Oc0RBaGyw9AViXhBCqOGdhyVHP/c2rUhv3cd+4vCHaT/JsFNfsxwQbjkQp/FBCOleJAHG9ue8dT
QNhZU17PMWYUvzLDpmYFMV5m9Mrp+Wtiu1FL7ujeP0NAYXvBYk1RLQtvqgYVnjfnDFo71WTA7QmA
ugX0q1Vb2ov/YyveXZYpR74IKGg6QqppZt2rcsTdOjo8Bs8tZuqQsAmV3lvWjINvh2gKTTZGpFWm
xw53WlimRhSa3PSWwnSS1n0REFWg5cbaM3QlTc/Rxno+JtQXN4jNxJoJFTZJp+cOnJROAIZO/0Tl
vyrH3med7uG4e+C4Sx6jx7KrAkrNiWsV5iXNFxokVHIRbeM9mo9GVBW4VftG41f0zr6SX6pgu2VG
yQVPQtnnpG/cXAyyFtREDGO6+MCaKsb2hEtVPxS2UV+0F7qaJG6Hw73GH7Qa6j3XTQ4KxZ/OqEYu
zvVPaqXTsO8IXy65wTRJ5lKZAmZz0JrJuPCxL9SAlKFu/ExUKD8JSIuWJV/g8N+ggF/hPge3c7Aq
UklqMhXO3SMGtdWZnPmkmeV0E5KgzTVw/OHDVdZd0z790jm1/zHQzuiAnRcZ2Xmik6vcCnuo31pI
VqFVVTjRCiYaUD1Jyce97YdNZ3/TokY1cVKmQoB901Xo8/atpMrqWHnUe7sRp768PbxSnOhKu933
Kjb99zA8Jh3g/ucRp7r/4kF7q+mJvI0fvuFVEmgA9Np/QlCdS8/xpEh3tVbR6qZkqw3YcXXjUVNu
T0F0bUWG3rixL3p6VIATpQLENfZxW0496tEbRugRRRW7JzttPFiCHkX1++04KfKOKCySvjHyla5f
VLPT1GjiJcPDAhuGQvBrbhdv3rA1ShJsEqryiqYVBWlZaoL9CtAvCYbI+subTV57+KZ9uc9VV/KJ
VA9Q+sGisxIFnysvxjhqibT5YdkSQyaYi3o4u2F7vduD44kwv8plhQoTd0I4McbgJ05aXoW5ahAy
nfzbbsN1LU2ucbUqI66KmuDhPvnOIAHEaZ4rwaZUVvjDlnvlxhBoG4U2jSzno9dAyDt8y26M/pAC
BGz28TzJxpnajz0LeCnnXpff7nnuGtT5gk6+GbJ1moOGMN1zEm48zhk5lRKiZZAO31H7mHHHPF8V
62dUXTBeR/Sj0U1eDll2+QBcA4D+SxGgLWv4vRCwiGoeeJj+7T41fNxj637LTcYANygjxgGe9OkM
cYGMekPBK4hjezd9xPe1bSZrSe8HUNzt6mE74u8ZGLojyLfh0aGFqdmPfzEoaiFhdbW1kp92CFE4
2CeboVmw4g/a6z7tlto8OANPsmrOCIOUOuRrTNnKfU5+x8gL9TtDz2BSdWhvI/ExpEBS2zZ05DKy
OrqcnK/Bi6++68TQo+wSNTgNnjDSRQQBY0var9sGC0QQQPXQmFuTwBjO0Cx9OJpeHgQKM6Aazo1g
ukmG3oWKGA621vaJDDciKvejAERMFKwwxhuHGLcPq1oU2yU8iGjR67ZWK7JjX5PUAR1sOtbZ6Jz6
He5+5EmHkJwkBywag24sdQrrZhJYeF611xf9ApsKi/tJ7y8z67EG3sC0s/B04RY+aclWunkA7gqB
6ezWveIc319wMCQjCdsVzZIQzM6rbZAt6+8dXimjEbGewkecAGeG+IJFsiXvZV8/gO59lYsV2U7J
wocMuX+vNq1n/MSwn6F4YAVf0esaTJpcKHTpBNrBzBEG6x+hCR8uT02zkGLu8yTLtjSztWLfMkhD
tNEv9VFKisNsrCnd+UULQscxp0id8FiHPrewDy7hBm5Ni54ZZMbzjRsxU0uMHW9RFU+eDbhcmw2o
ytlJ6CbOGj4cKyfxfYDiGY5xqp1U0Tp4DlBQWbUjcKGfBmN4KxEFdQB7yRTIB6NFLNzz87q9Mwcx
4LzJ+hmJkqjCbo0onChKwOqk107KgQm9JEH7vHtoZwjOXdEAeSZTLPJJtaWm9IxTm3DnK8W2bZPE
h9IwZjRB2KLRB+PWqivE4Y1LuREZDx6G2lVpcPkgwgCGx6OdqK7DkH4FCYc+9uVkbXYDdvUU64sy
k7iH1ZMHUa6AVAtUT7CQTgbTgcEm4r5ZH1StBbuStzz4JLMK0dbM5MOGWkzXRgevRBiyTNPijanG
a618I2FDyhzOA0Xu4CFf0oEE3roPwMKy2LVsUvpgLYOXcTcntVWYB2lZRB0sF11kUDxQO765I/Bo
C+g0BUWFXdWa8LeEw4O999x71D86D5oceqM5MG4E0NrA7vdY1Gu0cg0g9KaOEjJAbxCzzKff9vRf
R3U5ivgQ0CIsQveG2ln0RhxCudxLXb2CvJWjEyQrbNav5bZ6SQL3ly4wbecuze25mWxuCsoLtg62
G+DaXaOLgcH83IS8dwhwJKM+S3ceBdz5OINgEFRONwnAhebuNQgB1dj8Trt38UvWb/71RD/clVus
UF9mRs/nFclre3AAJe0rd51hOW6Ln4vROL4r2KZrTH4nQ6/NF6ot/C6U4oKdDiYo0MNdhL1w72ZB
SZVnwlFkpN5/uRguipktoCDjtnXlmdHygEwBaJbdp7Z86jvMDJteRWW3Vrs54oegkaxSPSMXy+oq
LNj3hQ4d73xGhbGxfQIYVKKKpyVRF6gU1I+vlVKttS67laEhb5iJ9j+Jx0r9v90GxiemFv0M3wax
EXP+7tn5EX10YjWBUgsUaq7gI3F4lDpDu35A5SbgYRcQfIklji3GI6xhj5OURIJ7vZj6b5GOGn7j
DgMQYlWbc569BtpzpHiHpXMZXEAPkr6HDe+J/648tzOcDrVCVpDT+ciNxzK+5N1HSxRKw9JQIzoM
0cz41GZ1HwIbTvOGTv0rowQrln9EpT8ot1rsNjl2kmzJVzwhFhh3ca3z1+CTGiQeK/3SxdMGR32g
sZzu+tiAaUkm0aO0EieH7kQEWKhvZj+JtpuwX5TE3AtQnO0FZejNRTdBYzi0ziVNlLJ8M15p413c
N8zOY+EqhZ6JzEtfquqXg3W85YByYwtIxqnm5w/ZLxOboDlS+SQbepLFZOJskQpzIkgSybWSfrAX
SlQb/SlC2RgGJ3yg/bJ3osi0P665pUco+WpEf1BPbKyDcfSnZ1zEqFSvhzBu7m+y2tI8hlp0+T38
GRRDfOUnitZpQfAEJvEy1WAmEsPMyHPLpVrBlYvzEzrgmRCb6c5HnvGRyBuVFe7zrhF8le4C2Aqn
k3tIyRxojbQhxxhYaEksXkQfzZSn7wMPgEm6iuRfHnPy8Wv4w0tAVpfW0acGujfAOV8D1ShfbI2N
4PU88S04cbQMvcCs4F751meXuIK65uNneXJZXcp1+TYcbpUOdl05xVqnCz4fpwJH7FrEnLVwuCsq
FhEO4whBq3/GuIgXelmuHFVVLBIWpUa9W3buESP0BMpX16OQshk3kiNr848EHgaODRgc5T9Ps/Ys
WvSb7rmwXszyPbkYJ53IE/omoZYLB1CypoUs68sUT8uhKnP3E2licb0QDmkRyaMLV+97D3QkELok
NN/HRa6t3vY7hwetiMT/hpKBQJaFE20t7WIJuzB0cJgAXxBIDoYFKqaNajarxl9Kbzc1Tr22fdYt
kUuhv3MwUyYtO+PlihdYOgRkcRolXSE4HkHb0LzBFgR3n8cnCkF6bnEPBYIyvKFy05e2A7hI8R+U
62ZmDQiGcr78kSQiIe/88mPzjuqBp1do5e0qzvcGy5tNa16ULoqi3+077m2v835B7bNjEG7Dr2DL
QcrnnTDAZJSo8n/s+0dl1fCyqBPjfEX4URtgl4FCWcRKAzDss5KTA23Ra1cnRJQQFPEE6idgZ95v
Z7jSN19UAtgIYYV7QzxUS/rLrt81MgkmIsFcONHY7JzWbWkDhf6VQNwDUuBMzP+gc8DL5jyXUhhM
9A0XkJE/H/ri6ono4SxmGs7eb+UUajiJ4raoG2ShNjp9dZFakQaZFEbYbuqshZa8n1BPUSPGtbaY
W2TknQzo1kLysQK+DvT2YnhPpTwgN6W3DeyoZ6M3m343VfGZgJ8CojgHX0XKuci4uLmOaQyTIfQT
G2fAnfI+5jXTxOoZMk8JTzolLS/VunaJzLXofchp8hCdGxaOfhHbXQW9vwSExzh2h+/TZICxE5oh
Sfz1nQfPLuOm2s7yrfhJDkbFaETLTioRta4CroL99go+bnKt5BcYPyMf01WhCBXc1d6zUuOH4KyN
ZKgNqyJ+a8OlYyP9wytFQrJOrdzQjg+BLHsLn5g/ybvNJloKn6HLg85X5L5XSk5Myr+3u5R8tSTy
RPXIaDz2IYcnGenxZ3M4SzJN+z49D37aOl/0ByMc3TZv3Ac4NxCoQHESL8UNnXqw2GH7YaNFpEQf
3AbIsIKQsx3rRMazAT0wPz5RdF+KasuxQoPzwYl3gvP0igf8PlF2HUvo9Lvh16NldJTEAbgMxfsm
46n76ijiZ+YcbHxXFxMwso5pheROgk/5uWIfUPYgvo8J6SU4aYIcbUzTwQ0Zapt5MlDc6i2bwhPk
eP8XRnWFP+RpJkYRd9i5HyJj5/Wv6nypnbCsfoKPC13muquWnYcpR8PeGwipLkMve4AtbT+Kvsg9
QwyH1gh29gqc8lyXYZbI17Doi/b9VP6Jeig6CKuuwu+PID49Q0x2WdFownqQGlcoeYchhLG0rcYB
mjF5ZUAovF5hCz/JAuhqT5CXT07xHfYtxImtcOWFT8feNFLrh7EtD37UX0t/G+CCZBd4VKi17vyw
A9eYPuiCzRmEkwT59vPgl6MydP2uMBt2VfsO8sb544KIeyxGKlehqxEaFbDE5l6lms+EMqjMiq28
SVJFVNVCzwy6X0KlEaHzMpq8wypGLN2xk78tH61USfyifPkjaoxHYRDWO28ojtPg9OC1FozhhUKK
IQZSC8EuxO/9AGdZAsT1W3BKVkOcJ7IdXRl0Qin4RkoZJNWkQoGIrrPSj2AO/rh1QcOPqfYQeSuj
T0UI4YnpfvfV48TE7bA+fwRW24ic6wSZ3RD8DUOuB8Eb2mUMqy2pM+N2vxpfdt7xJ4cLba3SVWSD
BUC07kzcSbRn0Zz2eIsH1ZA1iy4o3cHdIayFTNZLyPZqyfplGPl2pigdHDVobaWJj5Zk9b+FwDj2
7Ljs864cy8/SYwEUkvB+dnfyDN7bIgSrQJ/YLZV40H0o4nBiWOocH6+5O6eoL98pBa05P5nR+8UC
sT15Wu9hamGsWHXOTzzrZ2zzeReT2rfZpwZkDPbKecYchl9OfKDl6pnqAuL8Aftze5uQdyP2GwWY
y2AoXvOyk/o/1yfOmvP2wGJ+5YmQ7iZC1dDBHLnD/t72N+Br6CFlka3zF0bZyRNi5FpKZT68FqVK
4qrTTnCfSyPgC3ZH0Bj42A3e2PPhUi3JHMNYsBe27JL+jaA7hJfEoR1hqlUi6fRNaJaG+J6gRhjR
BoJx/O1RmmWyYKZc5IzXUwuWvzKLHJJBC9Ib+9ClGqZVJd8Zh8NCbULJr5R/G4G/3Tsuzt22uzwl
kz58vk4V4Z8dznoxmCC8S2RMmbUVfAZp7AcB8SziWRQscEXgAm8/EkZKn7bYFbnudlx0jBVx/WaS
+i0lBoIbJMMs09yvBS5vO95FT7M3LRBR0eawjey6sxvy6cqF3unbQx8zlW5Iy/9jmswPPdKNGOQ9
UNSqSXvBOqmNwBoXSZ9cF8wl7rVv2bPp6NtF6nlia0esO/KZOnqu767NQ6IPPNynMMTQcpjjFeN7
ngvtuheVVdnKyfXvz6ApmMOqmu0YL29MBmx+e5N0Wojem/0b1xtBrIh2dxP+F6q9avukjUtvA9oe
78bZDjuB7nMjd4YwjGx7TNl2NHwhxhxygTAooUdpfsBMp7yZQiYBjdIEDrSjDbAa7cViAjvAjDRY
sQidCyEK8VgatTjaYlXlg3xTdL3k5e5K+3oQzjwEplOue0fHmIxeP8jUt2daP76cXTavKjTtzQ9p
Y6d7xXP7AGgow5y8TvjSIVxiUCA1w397UNOrm1+MMFQu/+CPLgni1AY0IyuQT0rMq1S30Iz3kiMl
ixEPi3sCjewslp1n8bLODlo1U3+N/yChxRAOU5/u9yWIyXRUdeZuZinWO5y2Ytq6JxlpmOteyNtb
QvX2cZVMGLSsydEU0whucq3Ndz5EJtO7OUV0eolGxPLr073pJEJoyxBhkNAUFK2FSJyNZ/vw1a4M
0aNj68L4ugZYI2DPPjHpteI2o8ozsRc7XUvOYKa4o8McjY/vPRzXiVJb11HEcypPQPY8gQIbc3HH
DmfBIfEJJc+S7K/oMO61zt/S0JQ/7gbfqJmwV/spjvIr2O20K1i/+JDPI9B980a7zXCLQWTSWgl5
jAI5WIQrIJQS7Ag+Lyl16umWZ6B1ZKcTQnF0ITgJoeysmTgpujpSX8o0w28meWGqnLGbc7/JuQhp
ldrtnTMmAhN39pTgT7sdJSEcvMoG9qkUighFY4/9xVo4o4n+tY9zdCbAGs9Z9QEaarLslgvlM71h
7/P27CdlZvpiCi2wkP7/EK1o0chbxARGwDPd5Kj1iRYxvTcjN+dupG3uiwtlSqRmRGtaq88PePOm
X6LkpKPkFrvWfGJ5S6TAq3RFlsRIvWQqjmJPHOOnbQOIMBLrJ6pJZEwZXf9KsudTmQ7obd4A+/FP
IGRx9HYegUoPAqjU4EXYRHppKk0yuv1odwve/SSK2fEGr1BavGfBcYXicAX7TciOKfU7A9/XtQkJ
6M8KpRXqNsmx+RKv9aZu80oUo//wkkyuEf0SviyojCHxpW8tXtgw45bFRefCSecvX5QbMscjC1t2
v7Eg/BTvVKsStuUh0w/2pdh/3RFJuGFRx2e3gVpc74RSCLoelfFa14sj+VULbwRPs7A0xAqx65eA
9bLOA9cBH0Bezba8Z0Qnjsy1ioJj7juQ7Zr1wxxalvvuJNRlxDq9N22Nq1kfTI8cIN/gX7rXFWEB
URohhpX/Rl06xNdYwRtmSN8EA33HT9P+wHEX0pIBlf4XfpYllKfnKGBOpjdY0z3vIXyifnHnZekS
UHtFSB0A1Sfo+MmZJBCMiRHJ/vfEPJm0EeyD8gDDD7YaQY867cYy1Uzq9RRtXvyJfQwvszlxdQbx
7TVUofHY+joxbaSU1Q0ag5AtG/Y/vaLMyR4RcnY3K7lv2wPBEcBT7eJac8ktHXpy5QyNNI32WM+X
6jtqR6ixsGSYjJM7zRx90G8RcgjlybYtEFfpW5meyoxnQCsUxtMcyidK7VTmkkp1tABrVj0vMWuq
L5QcBoVB/6ckxrMkc97ipSoqPV08aRN7KJ05pnleqaQ70vT1VTVGBp7sj7R3Opo2i2kiusjQ/c6c
80jhHZMTACXi0yQ8/juyCHdJG6XBa+l3LaEbkQwOXD+BmDShUpUbNOV6XDFM+mfLwSbiSISp0us+
a6/ALm12uZK8GtUIpdVHIjJAoHScCzOtBIY05wJjYAqM3CQZ+JrrjtfRq3TowzP+jjLH/k2xPVRv
fPKIBcIGpIRDsdIFLixCBMI3mNAZ91RyrhdqcOezMRjFBIIj1AWXw5+aKwcCzqSUVn2YSz25/4pD
lFG+26cx2UFxNHSqGNgFMKvduos9r9+Gf2DUSKJ/SQkIM33Tcp8xPpTcolzfzWtIo/d6++MEBt58
vuvpaXGcfWMsi7oiCjGOOymliQ8oOCXJiAAoUiXxECI7Y5bSFSEGLMSllJ7SsPlqSf6rTp+06cGr
3QaDaoEfQif71NJibpttC5iwwuWvgrz60dRN18k+eN2h0QJ7dRwHAy3DawdA2MowL4D2LP+jy4pK
3WnXowtQoOI3Nx87QebSmHXnnaxGXvxntB6XlzYDQ3PxbsiQY4JKJzmzj1vVufEV/RWOMbdJLgkU
Z+st8ra+RrXTcDzsYmlgGP7p2AEb1JGvclK1Iia7O3fDDvY9NCz/suH4lCbSlqLJWbe2RvS+biaD
65OAZ7zn4n8uqbWDvtP/ed5FKWlcta9jHfYLMpAFFAsgH2MBeU36CVzX9LoWMIK/leTS8pdinkQu
BDtKiPa1uWrV9lIrYnVsVd6vt85wMiBMJ6kVtj7tm4LZuFiRVsn0bO1MKOLIgX+dCWy+1svflWnl
vYd5TnlHWbLvdlXV9ysrSuTwglNQLBNotwR/7+Kzs9tzjNzgyXajxNF8JrQTkq33KzbPOJwM4Atp
CFrLYQ8ZojHsEv/q3//LezCsbqlH5KlzY5xztfwntJ9OnxYSMuL9ad/ys7rZb4RqIkz2hjZkAPLz
dhvL51SWur4GCQR3DPYgBj8qQwngAVfocfu+BUeUxyOXm4EY9D62UEHmeWP/Ajn3s4Z6kl18VM7a
MZSMI/F1jOcqLM9JYEyjeMWFw6DiKXTtgoMCOS7HITxnunG6ii3sWBa74R1OtZ9k6PLV4nwS9lBA
C/gctVgFusnsUmlk6/Me+XvpLQdvN0Qawif5j2l9P8+j69pfwYfYUnWEyhlAdkG1qcq6O8P+UPMy
02MxzKcCfwylYsoUxTBfFuZjXLwT7WHPUBrAZZ8Zy7JTgHhGeDyFoNw1GSa8Ovko6WKJRkcSpabJ
pOyXHTbQDnJUH8vxHGosDONj7WA1WUZCFNS1WylBMFfyKeXoxwpS/YKxuvsZoaCP6GzE8EKx0xu9
+7byfc/83dzh4T0VHVu815HDr+blyKxr1nbQiAK0+TDU8N8BwxbK/hVKRMyI5PBKS6hx1fJygt0p
9jO+bTBWScWVeHbeea8k4mgU5rfrpSVOHaBAiL+RBmIR38ZOs2dNQ8dEglEJc1rWWqYX/Oy9D9vI
S5EqZu5MLkFz6fyGnKA4MxC84rYHIVmNO3PYqIFkeVFV1eXKCchKty1K5VyzrDOYi7t8ueQtS6l4
6BKGXgITOBNv6tjIEXXr7mFZNDwG5FiQUWsc1oTLixyYApo/edugwuVju0MhZrLX0IJayeA1irzj
60SFGBUepRiQKYmfwnHOMLtWrP5pT3141Y1ygK6tm/lpaPmzyJO9ch4u/nXih007a6x8oIy7IZrR
CzWsT5VIQXzUA5khqbcZMr2MWKtf/UyGsUwqUkBi4CPlgjNHtRU1/duKnK75bd5YJJPtUsyxOFdI
r08zc8Mstu7NK6ifKcpXid5hKXF2SqJqaxVVjul8ImFaZ/+cZHyb39vp/UHL5Cqb8VUvVkhV8gYx
2WLE8r2W6NcxO94jPIKjtZ4TzTr3SQa0EoVEuY/8qvTDXvoLmE8MBrBwk6+uvJFwPMDTYK8F+HfG
ka230B39Fx7DgVVyFFK683srylYzFGZH0qx5PBZARFbdvZeB7SD6eOvMC2maasDStNibPVshwlR6
U6uFlEMwC88bURfy66GFjtoTOZri5GgWSRKFHHoVpSNJ2Yhi1LzAO/lN/m+DTa6tR6izWuZ7k42b
16wutpPt6HlCZfS+05NLV+ZePVFNrB8FYtWegALb3hzROnqPalehVZK5sm0cXgnuDa2LgtKfr99U
CePT/0gvkpd23NVLXckidt7aUUjR94Hefy2ygoMPD6Ewbe6WHNhQaOrUxoteUGmV65qnz7J4+JVw
w26P0XLDQTwnPAa2/ZPOEBiIqzT6pkCvqTRQ4cERAp3NsLxKDtM84CXUh1klL/gzp50il2VzYDCc
e3yCHA6QaRa/UIdpbJ3xF4dRkQVlsRw91BUKMHFrLLdGOt7v3eWDLB5leRk6VDZZlx8Redrhs7j7
aGBIn/gAoFBQCUJkWS63olbzGdftzyTuu+aOyRco1rgftUa5hkkn5g3wgVLtBGBNsBRHSA90Io+3
WysR+/lcOZTcejumiKbGuxMWf1nay6a8PmKOIqOLjs5PHVOoU4vOvL0uoExdk1p//Q1pvX8WCPN2
SooQ08VUl45tuQMsSG+VldCOfWL+9JQyYfrekMz/zS66btBwr8nWftLC/QwQv7DyZh+PdBTgWvOh
ZxEKZH8oSNBFQnQXxJJkw059Bww+coFXgFyX1u340RkmIngrH8qO/xoILw4nwOGLTYEss1NfPEg7
Uaoc1ugg8sIIiVpBA1codPsdBFUxbkWmMG9tkbIvnnGNku6r3WBCTEuMlXTlFny5+//4b5k2vHPg
J98GjFQIjznKyAWu+on64ZBDN6QWWpn6pQNMVMOMRcAF67ri2A7nsmKt/xGOQwaNXW69VfnablPX
6gc3BhQ4rKoOWO9SKDfuWsoGLpNFr+YEJYU8yNZSqX6mRimqXxLT1VSa70GwbM2VhVRi3s2Gw23j
zSJF4c8Rys7ri8nQZwqDcNrB3RrtaBKsiG8fAcGu5661Tb5aKZxEA1K3UHrcCAWDg7XTncONm17i
f+7opB9ysCIJX+y61Q3XFXTX2HtruCZqe4t5hMs1Cb+Cv8zYYdNRtZTOzpTWgxHkgwhxm3ghVWIe
VyV4U3ZjUIWWpi2ktmEIGcmS1WlOMoUpESgXX0R7FP/NJg8llEo1tQxOBKyGn+J4MirRYwEQ4gcT
BNb1c1qxJJz5zmMt1KPkF9bYAvPpJkJgEmpmG5WtdB/y+VxrdXY94zL/0FRERyR7JoyeZcQlmj2E
HF3SuQU+dJMGyKel/d4a7jSW4Rn6WEzuZI+Va+TCrqVjoFkUNSC3R35posiH/fRhYZiqm+mOHxcy
MbkhX6tHkcmqkV3tpu9RexVpHtluiwOJ0ijHWela9bZD4sl58z+LYi3CTcLFu+YD/7UwiT53ihQn
yeLFTYgjeuAIe59ZzaOlFTX6sTZKhs+TCRZ+xg0I58+zn0v1UA00ZqYeae/VLBjpHEA0Ee07ovPo
NRdV7UIzZ+90uOoJXDYKHJ3nItnOP5Yzcnu7IDH/CALxVcT8mr00TY4xsPNBxwRG/+xhoD/0745b
T7j4eDqaS/p218ABNWo8+BYKw0wqZ++5/vjMNpfbrhgFVCnSGp1EJyGFge1Izt0OXVvjb0dSvNa1
KNM6+gCqJw3w5IUHOVn0X4oGIL0SqsGJUGLNX8Rxk1EpDP6TpyTcX2aCaciF6s37XBgWXwlR3lu9
Zj+XL8FILPCG416riTwUwFFMC1GV4ApfxEPatA+YJF5dxyutNWM4o7HcVGA/YM7L8MacpORlRr2V
8kQ0IvJij0omisb2Zt4RIopqgJCMQh1xeLFjewBoRlJkGyXQb75Eputda9IhIBM+ZqQ3i60JAOVs
CPOHUf0UHRmtgLWtLYyEXg+n3C0OhO7ZlrpB/RAWhMSZAZ79Bz2onIfkiy5w9jidLcXdbQQ2LpV3
fxK5bUux6CLaCvIQZMx28GDJU5u1M9UKIrg02NVzhlmuDfxleTwkgSoMeQPlcF2dLCSS7aX2Te4a
bmgwDDQTvsIHh3vnixX1U4TZbT8PiGWJOasVgrSGqSSbsJcViMfB7X1ZFYOf7cTGVMZIY41OwEGK
r85CmeRvW21CTJM231ZhAuk1eR0heg85TCCqFRU5GpFJlhuKC+XcEULChnQlad9zPrD1RaAgKnu9
FtJEpJc/EFIRjjcqekdSLi6OyXXTFM9DM0cwRHLLcqGiQxexAawHpS80sGAH8lJa43eVBqwWnV0S
Wsd4BzJ9PxInkuFK8E/hqbL/To9jF7Qg3VCzN0Z4CoSE3rSmtAh1okje6ZPs0rxa0CQJazUFexP3
fA8IpQnYaOewROMlJzF2zoN3MlNVYN6tTw60xuaydipSmWDtQPcQ6Fj/14je04+aAxSVMM3+XSLz
Yu1LiWFoK6S/toQNzHQf+FQk7jP391J62/V0vMUNcsKsn9z3ZrHSQme5Q+mhBrYCWxH+m1IEJ2BZ
0p/kD1VUjfePCmOEwp2hYicwtHuB2Vjk/SODr8winpfgg2p7coek1uS6LOjBkbnx1BiAR+f6Q/lw
keOmfImDcDoHPn6v6hdj0OWvtil5uX/Sav0vQTuS+t83GnQVWuEFZaWNHA5R0AeqFlT8rS7aIRC+
b9QXDxj5BuA0PRD1vvUGYp8uW9nQTmbbbypchuupndv1+3q5RxQzlEjuAnod2LV3JbURw/IS21Lw
slihMavpUiBVHdOQ/Mi0zEJrXE/EKcQC5U19B/75ZkFZXPPf40pMGp/teOmIl4gPu8/hobPkQ1fI
2bQ9mPIOe0FM3sof1S1lJ1rYJsySgQKi2QLd3y11pL6S3aq5NT+Pc5kzwMfQUe+6siVNiqifAc+r
LvlYZr0CJbhdZ9tsHkkWyb5RmDwCtlDrInxERrcB7S3pb04Go5COk8WChz98YSBivqudbTuELo/L
41pinEQIaUHZ6rh3PT7TlA7DC0MlKAzgNjK7d+t0Zt0IWnk6W0wkXZlER/cmVQ+rqnf4E6v2Qi7F
EHcPoKQs3h6NsUkrnpSwEJC7oCfK1msxhhLFUoY9brOZJ+O6rYqTU9WPcO4LLtmZprIandkwoYzO
7RLc3QgIOn6oS59ZOBXJ+Ck/hfGGBQs8Ry5IadbNm+upglmrPzsCQ7SFnQjd8IKWAECCYMUD+/QO
OfdkBZ21zjHMJIJ8doxd1CK6MB4tYKaa8UMsAI8e9sNueXQx9+gNNbhdISmmNzD9CKtcMPJddzk/
Ava6uhcfSBeG2/WMm4yTGsuFSftKHYWs2yX03DzjdrU+qs76Gkr+EYL2sNO78/5oJinvhvtS/v4e
fsOrA4IHSGffkYPNPgu2DGtJ7RnJycnnN0LzNLgndcHR5QkuWxUUtMh/8cOUTtPGRH3ZAJ+jtA40
xFlxZ4MygsLwBXiuWWpJf2Eu5wbiGIEd+KIwQ/pW0sInerMfARWDCKMjDGWCLlZzdqrvuN1jhgR/
yOuyrVXdBbzcgBR0L4i7jqH03k2Dw6/7mtEzvsxLcffzdjpbfBcW05sc+ahBfc/tS2pTrnxYlRDc
vd9JQZN7z4gN6vVv8re53dELeGeIOx5XaOenqWl1zTsm0ybA/zmvOKeO+2EJHxE2HYyxFyLVpdRQ
4KoRafEY/XrFJL0GUZH9yUoPe5y9KayMBh3wPomOZnL1CiodHOnvuiitIwsoh5RUJOts6YmSJjGX
C4gAGi9dHjbgZ3wpNXa4zob1STfBSWp+ZBokPsnSbQwQ4TCFhf8YcMaWhbXiGt1r86PdZKo7nxhK
2j/2mw/q+U5fC5W3Azsboq5Gck434zVlUMS6wu5gwlFrrtT1jy8puWCgi2t8bCC1zLyweYz9ll6W
hljhbVRDKSG6sg8mXmUX/LFVvnz8oXPLfKr81zl4Q1YTfncDYeu3635Jhpe1uyZRu2wNm8noQ3dn
GYpRMBGJfIkmRgDSqia8EUdUARf4BJ96DR+fD45knMJrqEiei8BkZeehd+6MsD1HJdvtMsi3EjNb
apqDLE7WcxJVc7yLk/6cgoFOsK2+iN9lQGjGAtL0iKp8dP9UkJVHTW5cu/WDlWxYKiWsEXADo2jV
ZrUBepQkWwE8gZoI/HFs3vnFYIZvCIaG1A0o64A4U3eHFAHCyk69/Agb51t8TTE0hJJYWmxoJnMw
eDqizS2PjuJVXfGWvMVPaFM5vghfJ6puvbJ1eBGuu0J0wqLBRH+3RRSxent2wzEonOY5xfVXNDdz
bQ1Ru3Epv6U3TAM2Zd5cQDzDGIYqswooYIv9qWjaHSsfKLDqyDNx59E4W/efiNqDFARsF7ZeMgc/
x+pIJDR+s5UBG7hKf+L6rGjPmjp1eZRrCRTUm8+buvAoML9vY3Nx7oBVnFlV9VduWBtiaNSbi2zQ
Q6lFuFICol0hokjeiY+5B8ZLBYdSE1dRCJ65UuDGnWOtJdoLtXPFMUJI9d41HzGa9/pk85eWQGyL
m096HK4pMH0gGZ9DGcxAtiK4UbJ8WNDOki0gyEBKP5s/jwaO/hyEQ8R9Q9GIQMpjlU29CNaa/h2v
HhCpHEMijXIrm3UImOGLBKQr06wPOSjQb+i7Nfw91qtf+PJm0BAZKKwWyPMGivZlVrUhDmnCoq7n
c9951+EUtYVyn+VvBpyEuR4WlY7yc7Jwhz4COnzdao92aJnRNgDQc0RlgRdYKerQ+Xf35TWrU40I
Rsjg4+0raHzJ8wEqWYKuDQYcYnMoAOBQrHUxSV8+oK1pzui+PrLFmQPuyU9QORgBXGh9YGJXlW4M
i7TXwJ2tmhyKyNK4QjwaV0k0zlCvG8jTgMUnzQ/pEb35uLFG3xZ02I1tFsZ6KiW7U+B3PxCrghFj
WYJ0V5QbGQuLZnxj7HeXJesCGd28FatR+CcP1jJSJvgmxOJ/0sYnnlI7LSpzVwRBQYEv3vx5pgUn
NXxG7WteOhoXfn99RLFD7EeEfAFPPi97MkMrpwdrDovs9tx3pMKtCeSo/Y1GzJ8PD7D5SvUHdxQ4
bYzr2aQSstvF8E0jpi+9uExj9xIm3Z7iHtsQbc7kkuD3Q3uzQ+eYZlUxcYaMk6lBNhDhfRCKTPLg
bKfzHJ4xw+v//l6zWEPMhYYZZ9MKOGCEgHPasUfGf5sqESv4YTZAjqhOqm1BUh/GwF/Gz6b4Zmz1
cHLeNX/ai1lCR9lpxwj60EAxwgdA++yBYudedrVm9t7m8q+dRLhva/rqnKj0Ro+d0HMeseFyyiRV
OyFys8B0nlBzPSjbXm0Fw6lF0cl5VD3E2HnBGSoxloutakRiJGJiNRWrGcrlVDJ5BZWAp6GtwB3c
0oSM35No2C7Ce7gMFjCSxUqxHzWgCeuRTJ4vp7YwIctiVhfyJXyZSswsm4bKaEKAFxFG6pjfo8FM
dU6q7Lry1XIP+M4fHFirY+QDFYYgm/BUGSaq0Lr0zSbv+XdpmM3T1TWvrN1Yv/TYWK3rkunWNcaA
J8fYW1DMW5QsgPeK+fSsuYza1DIyKDFFCbggn1e4Fb+evOFzU7Zwsqq2UosDzHGrcM7c0HW53AfZ
FwxWRBM/8UkGvMI0IGyIU9ze+l6lvTwhIJNxRh3YTcHy0uJ03ZUJtoHoTeQCzGGDny5N/ZEVkTJR
GD8tIrXZjKromyjy3AeiJVPG3VZpasGmdjDJxwKgw8q1Pf2L8cDEJ1cAbYo1TkbdeNKc39yZMKhx
cZwuHP71+/R2yfVJ/UNH4TBBk8wV9F7qFWy1IkMxWbTrClZGpFUTxaPCodjopvS6FvbeCbLL+6sy
sn2onQETMFJeckYIN6BDzM7zneKbrIi/y1YpvXF4fHR7Zeaj9uMho8W5wE1Js+yf2DOGloDd4GVG
csSeAm+EvQSZe5rZo/DULMvJ3cTGUTQRl1X3iJ79KrjCrY9Fa+o6zfuU7NPfUj4vPpVf7TZyIoSF
j//zz50DW09Uk0SqZ9xwC4lEef1kNyCir8tyMrOBiiVbPrcIVY99mPFor3U1wMPSAduPnRqg9j0I
67HPwfK+lAuF96dTVljRREdLq1UkueqoGhpP50rCsaPKCRMUak8FdJXmuSrlR5OUDgmPOIwCbJIx
NFXsRU58Vb0cHJfC4ZJONIabtqxD7ghLpsvxqFuALe71P4Rnl28LyVltTKjTS47M7mbQZOEgPH9a
hPTl2YwcZeVUVjM9llXvRe0bSLuawns6uhGHsi4wdlk5SLxUhPvw7+KUGMIHsFXDVmbjLVRzLCmd
IcAval4HQggf0b3I9iO6EMKRB3/B/LbScIRbvdvpSMR6k0e8ge8ESBz4yt1atAvI7X9r9N+QK8m7
LqTkztXSDGkwQYaYIFXEML6r17K0aq/BuOYZ3/SRwtb0NarV+c9IFuXS53nzjl8kWdFsQRIVM85g
yftPq1tK0m2uCdAWi8vEaUGD+3rx25HEEtX1MREhF1i0669RCRTAcOcdXbbAkGg67TXfqZ+vuCm4
KBzpnq21h0sz0stA6pk8ljc6vuhFQKl9jFq0tEOaWlixR1rgqtq1kB1p78LzdruI778j7lwKFiav
9UB3KOHS37MWG1qpvblVZwjCjzo8ZsjYSdgcSD6Elt0i/I2CaGNYCpWvReTlJ8zViDJrsr5jM9Uc
hkKmctLMxKTNeQzHrZsJbAXUCYbaoklk4wBLl+tGdeV3SYxwOoxjqdEFJyIUAYdrHEkglWrRT0aV
OLtYrZy7FQHnxeSSiV9zRTiN9kRxFHh2L5V2GU+u232pKkGdA7G664yIm5moiWP1Bn3SyA+UGFqB
ywct8P+wSDffzeHIu0CGXJEr2fxRWWNUIWLT4upr+i8pYhFv9viymL439Nl4W/qE7ICcD6Wf3HY2
/HJa+5lans9O9VR3wibR+kAX1PgjGDqmOPAhxBNbnLIJYDR0+0DAPZlwW9OpvweQOLM9FiXufyGU
N0+dss82EzK16rbF1Lh2EpkOAUzn6aMKrsRc1w4eBHzdDUGXrX3u557d7C0DnFWZL0n3qpLYcMGk
1vnQ8oEbXxoreq0akiz+xmOZe29Z/KEdlrWjHwPs4wtPKgqv96dGWZgNx80O8Bfl48eOc9Zns4+U
smaw0vQxTZGpIIQ/hO739Dq5jnR/WhODyv6AfYwh5v2iT+jJ/zURiZTjQ5ixtnH3bIGaQB2Khv+s
HlEqFLih989Z4JrEzwB7qsgVHz6ByuF8M8YCnmQQB9Xqkd1/PhYe8qD23lU+DZfoJxz757ZPstwz
DXq0KXdI+tPBdGYHjjwTRdaVcWNdxSRqNiau8g2/WabDyvoClo3uZWso8ZC6wLoclt6mUzp7dId6
5wscBjO9RF6yR7jurGnpBxxNAJol7EzrOSNQoA2M1HWmXggvfxIxRM/brwaMGxD2RrNC5bPMI1Lv
z9egmQES7rd+074JKbXjeCmbLbgQyD8GyZf1bK8vTE5gFR4qBN/HGlEeL+FVs4uF/hXUijuLOuCk
hNfS6IOKnicRlo9gSqoXD4EjB5DafXlBLUWXif8atOE7zrerC1CRcqQeRnF4DygX8uwO32/eG5VP
qXQj2PqMy3at9aJK6HNS5JWmXhDLG782uiSES9sSpuvwGvxIoZoMo3OmGYhrb+EgvLjIDchxPCXS
mMQ07Tn1kr/19QCg9jEFOWAKNKAyylFU0i9eIRMwMvKlnSdx8B0GanYoxLNyhm20qysXTobnh19z
psvVinPnPKq7gJghKGbesuo9EPIECbqviIph3HwG9QuPLODrRBZvmHJvdGiuQTL1aNT9VY+XgHel
V1j+4GjgR8UdVSExp5PQlSFt7NZeymw6NX5cR+7SmPY6rOoTwy50PNginYmMzBM7WlQJhaK3CrxO
zVmARjBsg7X9WFtyjp0ZgrJP/JJU/XrlWlzbiL7KrGCm9vp1erpS9CFOJKB2inIDAv19TeapnypI
Wq3vk/KTu5xsnqH5Td45jPaa6ztzWV3zf3hZghezaYcMBp3srrgazfuUnxMb5oKyCGvjL26UoBsi
hazb9DKNvE1kwNufzUdL2Tk25RD86nq916oDOkRDTe82qXJEQwobOd51yKUfzrbGHoZqsXeUzAqi
FVaP3QZB695WRGJqUWPDKaDhVtacuIUuEqsnnRn44ZB/ztAzgMoKrxS+BnLSxYWwlXNv34jUBEk2
T4F0qxU+TahJezFiSGeol3Ephg+h7tiRLhQ0lbgljRFzXZQGLNbnjL5xVTy4ERml1G63mmieyMgi
aqVTM7hELEvNgdS/FOdB/AfEyGuX76qmZuHr9hjouxWKnjnzUYRPnOxJrULVAWZdggbVuSSZB7pX
eQgnx6ecahjAlLAbFHHgIjG2L2IGJjSfUEXnPxzvhQGxc3SkDpriokPCD4ijyuLsNvsD8pKNsXSx
7DXlkEdsWRAxJ2DWILk6J4+hZEukxk9IlFhzowUC9+UfWoxmUUc0DbkIJx6AXZ8aXWbnagWNeWmu
L9KcfrXN/dOoaanwGZVGXSWVtY/mTOtMSD/q9RH9DnSeomEBxXr7KsHlBU+5TKHqIy3PrbzMgaU8
cXlAAvOcuuji7MPGVwfneHNJE4zj1a4MX1Hkj90IzBp6qTBmvcWREbjAu+HPnZ4rGnZ0kJlq4GGa
9LkU5brgBlTKpqfROaZB8vmdCO+Vu2BcddUI1caljLgq6QKQUCbv8YhqJqQRcqZDxDF5Tb46aQB3
XmWOzgn0DEL5kYC5jwXNd56oGr5JHc8yFytZewHT4IsrMtfTTfxy7Kvkt2FajA36lNwXZN0EuGwA
0MoPYRY3BvHQ07xUEksCKrdn/reCssd7VaDoWSBF01ER77SA2cHd9OJXZL2I90GJXoTiVV1cXuJf
+U2yqomr+chF60D/7f/VKFM663ab0kNAhUhIaazzoI942ScQU65l8u5rLzrZ6KVH+icepc3HGF+7
ukmdtjJ5CXSh0HbLJDfwFoeFNFtN/RXlF/+0MT6QiABU8lf4cn3I5GmsmO0k7iJ0+NQxtLRjVA/v
FznHZXHZVQ7aKIG7nPvXViRswAKGnPvqTXLUGzsbeDrAvzAkug60l4jKoZxD/8hpeizib1r01ues
Yq8VVtj/ccEtIkNkVFinqJwkSHvCfUWVLj9TFqTqlYsDTKvViWUGQTmVLxNkh76TmeTOjsHJw4X/
59PqSDzMA4zHOaDCn77gTNyoE9UnvpoqEZg/NefAm9vN1/STMTOFYBDO6alkdQeCu2Uxg/VmsIQV
SmtAHcx0e+oVUnNsmylt+PQSqkl1PNuCgpdPxUcj5IF9BQ1+MfF/1pKVfd2WrIeSJgLEaVs2R/aT
dlEAKURm0286+8lyYQNmscv6I4oPMmlSQafyoWfVeM44PANxcExn6iEXhwSq6qic6MuJ9/8gvATc
zikLphtaqG6uJEZSM5XkK5oQYqvdXxObRXQOtNrhJPLrVwQL0o0/aDK+3LDIvaF75nsQ2p1Og1Pp
C4Ae87aY0BfjJn0RJq1Q/8piiyBQ/O5RYj1bo+P+jBZ1+bp5uZ2PrcFihBZoF2y2J4swROoggBK1
l2K85p6kgQscxRbVHWXokJhnavNOu9hDjUnJJzZ3FYYFlutsQJUKKQOmaRIxsS+4TPWJ4zsrWijg
Z7FPkLLapJdFuFLA07NiTMi6Bk8IwieKOyxCs4EZYM1iYDOwT4qha4EEnQcFhsedtGe+R+fVpLUm
LM+XlijD8Pd963+RTuIj++B5YHBmbh9kmJqXYTJ2Rj2FmIBmINl4yw4woEIkH4DkBcS3kaJQinC2
euT+6IAESDookjdLpS8ISVyiC9YgbzGzpcusHiCKrg0MD5jQP/18g1msdoLJ71QUw3jkP6wuvGAf
kbhHqgp3SXjqOeln0AR2253YuUUq20KddIFYzFPM7e3G0YPbhqYA2wDUnLLenffc8xy81loVBCt8
vExDIsfWZOhsGV8aAMvc/7QYrLnFLLSmz6w3+Jc399QS/nv77h5IGAhnCSN6i3ZNQTgYaKmy/w3M
4YZwHRm/GYWu61XvtcRo4ksYe8K3h3Bl91Cy8QSEb5zY1fLECfsPR7DRx5dGpM+ju1z+yhBx1R+p
BCPX6e9CLKd5k+4+L7wAMoD3VyLs0iJkrrFNzBK50bCffXs/MXRy6p28usmOuiUemYB0zmLtPiJK
9f8QltAZEdFOSorU/C9gczk/Ab57QyXq1EZIm3Vdk28tfZthbvSTtVhFBsxl3QzU8JP2JL4f8DDm
zz0VpRX4ymbta8XxKKP3q/lfzP6Qy74eTrnUvTvJv7Czie4vmtQalzV9+843Rhmi3sHJ7eqrg37H
IeECQVL/9RvRDSZnf52AsUicjf6J5wQXosbskoh8nExXf+hM+Y4r9NUKX6fHvfCZDI+BBG+Y7z0/
Mcilxz8DHHQp0+jTWaxVUSENQbjmukxCixguoY9hqV96cj8SPVregn27bOw4axustvze98mtIfVV
jKAIvCbUV5K+DeF2uogioJv7z75REdTJR+OD6GqoVI4pJVOVZSizcxlkPKHkK/Rd4KpJXKEdo5uS
pxJMamIGKzNL/Zp7hj1kDOAVy+PU/5b0ccQFWQpFPWHS+joiRA1xlM+BdU5xSfER1j1eXGLQhfs8
MT3YsaxbjtMu3afx5x3p9g3Yt9fuI8vOv6DS4PGM0zkt76nXiVYsCuPaqwh/eFQQMgh/Feitlal3
PLN76Q5xjAuvMrQG35FrYctGC1mrJMe+cWXf3iWKaSksuy98gz+Nm+DP9alkeGzhEorrwCKoJ9de
tTyqVOGs77nHSYVYicYNjdjly0+fymHURESSh9Mm2EXTaoSH11j2YcsZDUpFyg8oFBsNZMTXsCRo
+vCpPRMldlEL6aFfIfYzeoWt6e5mx8hgxtyZpEIREhsBsiIJ/nTwRxojNhDDGz1Nt8P8TsilH6h/
oVPJnxpx0fwRNsYpGybfCVj5JohuF075Rx7iM4v+MkNBsKu542ekTocLdgqR+FR3m+Iz9se5aJDm
6byRBA3yx2dJuGsZ7Rt/dgb1QojRVjFvIPCmiRlT4gVsDtf/t3A0kqjEAlLEobIifkenUMeuHi3O
ZmCCCU9urb/9Q/7OXhKMdrk9oFlbyCzb6RNIGwoE7stYjJlonc9EggoLSiYIKfruJ9bkDLvw8pjc
+8rc62/Z8GExxryYsXXPtW7hh3p7OjCtoOjM+mHaQt88YCW8dYjbNmEbRCZcUC90QWH+h0wqP83x
O1P5K0+ZIQG7DNUi7aAhJ7wwDA3SGEFsEbw779+OdsDLTnAl3OhxO9N+A0hHFHt15EBC9p1ONc1l
n5/ScNkOIF+FFMdqscZP3PwoJpB2fYdQH6UjVp4dFbKAFjyNVNZ0Linp3wdDjHjHqufm/GxajhKS
qPsykoqt0Md5AkDCTb2tF4dL16Hz018P26hy7LhGZZp6VQW+zVxwZeClY58Pn4LP5pG+sn3XrMgG
5VVhn7r0Uq3BWAr899CPAz0dU/jsN8lf4yJk5Mk/3OPNPTpwf8HhCpFgTp+DXXKrcl97lbZ6Oh8i
KWz4ngs+BTza81k1rr7GJLCFP7LUB0Hzj0rgJm2SNCYIrQVg2AabJ7WZ/awtLqG6XDkOkPrMPQhw
Tdktny/gtTNG7prkwcdhTPiBu+/y1edqgVSNB+qrZtSFwIsIuYSLDPO84Dm4KQD5RSWEAF+HzTUq
bBFu7YbtqdYrapVPfXmjSsDi6kbWMCv1cjhAEK6fxu604nDwq1S6yTOsY3gND7lgtp8iE4U+zuuT
zHaEtZjPfwMm4D0Mv3gXSXrsPsw2YWecx4ogWljap0NFtBY5aOe2fRaGHxLX3+aGvaMZVkN5qUoK
Yq36fc/GmDhhx3RidWZWc/fVUblc7F385NG72Dfs1sanrAhKY7U1C5Cp/WRoQmk7YJqsoubeuLYs
8uCgW1lwn0dcdfk4e0SDJRqLZz31ssq8NJNwSz4V5Q3IU6f+zmg85o7ebYnSUi6dvxzJa5RHgeXx
7n8GSgte7akbU3zhwBXurB5SaoZT0G05FL2aQSqfvvw95dUu4yoTsywPvp1hzJ4gsd13PU3YTjuE
K6ZEPmkqnI3z6uRchI1ZnYkN0zcTMVta+vzqBMNeG9T2xL5/sda8SGU2bEvOLKLrK6bP5bh7bdIp
/jALsWZdMmpaPYMvSKlQ76E0PhUdvMrZhw1st8Sf8UhR0pFJoUeAsVbHfMLCFJRUV/B9M5GsaeUb
UxPQ6f/4ot9sSSXv5WZeeh4/c0CHKzZ4C4TZPbbR0irFvuLqO8yMcArt1FGL/7XIP1hEGo81uk/f
8TjF0do1FTpMBjVqOaWpYt2fMzidI7IigMp3ygs4PYZysXIHm6MxSw+v0PDetgambqm4ro9YcJdr
Gcms07gUU31USeI3e6iNluk40OOZSbBq1Zv/FF0KIM1+oJb61DboSTFFjbcth6FeuRfWIieGryXU
P3eU4pmjUj4DoxIjMBSG60C3sqHJ+HMCkPwKIl9TpMnS3gMvyJouICsWmYsWPXUx9BY/QPv2r7lI
xf1RfPD0oYqIffUSZ4AMdzwBZsKwBO+4lDLsLzxsVFiNXe+8nZY2JPsdouDlVLwkgetEcF0jYC5w
fjNJV3JsipPgPF3uIoywvqV65LCXWlq6Z716jHdBPJjx6cM6KvW8LHAQdA8/lI8gzc277uIVOIcQ
bgnILB+f9kgjvI9bxL6UXUmphT5L8PHGPyEW6bJhwJ7RxTSlnnPPC3AzyXR/0XujDRObUmRKjNIp
ICZZaQwcDSCrDSvY5j/e63rCdJGIDGrl5w9hViO0f6OHOzcKnVItn8FsDSr/codrRz7CbXkEEOSZ
DKO1zMCbsfditQfhQIixX0A1DhdRreBPUCNOWunFwYdGuByOo2VjvePYDo2gvALhf9WfLwGjyOqB
gAgNG+Fmz+zDHBOssOUkH+V2dJNV8GGLQ6vBjq2ckh/JzZEBFmHou0Td93akOXqsGqSrN5m7wzeg
qPM810Ps82RihI9+7BF9+XnTl7mpPWBDiviVvlpMOgs7pVXFkMpxSNeBld5N0i61fSe+oIrxs/1m
ii3fzDFYa1ei8cbHSx5Zv14R+sAu+JYDeajVOjBg0qceUPBplPxnq5nRPkjryJuA8cN8BI5xzKQ4
SSa7BJpJRICUEZaYkfxjjX4HvXcGvzY9/6xoXyUz2vRko8/v/EWHHCFfQ+QtM4QxdT7kF70MBYUe
ry3QuXvVB809teVpfCKqo92/WLQkp84+3ZmR5dwIqjLf/HnjI9Ctj7FCzBEDDLMykYB/zghSEtjB
IxI6fxrdxnhJW+/nzgns+mPhaXQ1sAenVgqf0ktgO+/mqSm5DiL+Arnx7OoNgFjq2gr0rDHvrZgT
K5A/Osb9CSwOLBZ9x8jieV+ukVaUww5HUH/CoBQ0IwZUos5bb8ZYHkz1YKeEb4eCrj34ej8Aixa+
53lD/BNTvPIe84XYJElnFcNZHLkHZHMMwnLyIhZ/e3JrK+ZTfHeLQ1LSZAAPDMibbJ4kfKlF8Oft
sx/XVfxrrA3HZSZueUVnjPV1dc3CfFhLNLT17q0PVZ282np3XwX0oj84EmfvSm8w0/2O2XojsQAj
hB54I56l0ySkvZc3iQGzAYWoYbclTVBHKMErlzdBNncA2VsZFMHSoxMCqZQcfi1i7nKCSb4iG86b
w+3XJzR4fSvX2NcJuMDi2jSkLFGcDw9no3Z+jlYhYZ24HOyicPuin0YTtvNycFa7IQwlyMMpDu/H
ynQW4+qqSawtXaF59q2WXTfVo44b1xKkQrxfVdyf3QnYZMylsUE8uvtaw6aOnzgjlBZdaKW14HDz
8oF8qa7ptSmLVw9MDwsGiwLorYwu50gK/NGbIIJyFOidQLQlFExerzl9SYLiOEL2c8vH7ovy1/2p
cFpv4FrJHSQOKQmlwmEEz9Fs/LvDSv+nGHFg/Ot62Ey4GkEFb74A2Ef0S+YNyklfzYeIBcBAMuoK
SDzJwg3zRuSbzJ6yzc7YnXVbUn5hAKo47SLdksWa7ZXmHja44UwOKvUz0Jm6qAq8lulmPn1x1mRV
KyTfE14aEOz4wkYvGKB5Sz2u+Y9Ei2ndQPCNQAWA2lDIKCJfPcmOntgj1H2w9pwLZ15qaFx2mukT
e4H3cXWQ7BVwJBNopAvt5AVij5ev89A5m864ZaNUOclC2OQVd2SNdiEpMcfGzjbxAWt4hy4jAj+e
npKcKjTof6YzA02zL3LXcz1e1aQsuc7aDdakn4JcG4W3bJtW1p2dmiIV0M1kfsw1EGdGVPwW7TR2
Eni7GdaI5TVnk2k0HrKR6CDMMb6Kukj1YUlryC01PWPLS8jmPPiWX0h7e/RTpx+i6qdgTKEiMcQe
KuP8WPv7EPE7U82juxa/HHQaOOPx0dOh8g9fRb4n3CjYBVzd3p1oS5SXysdCnccoIyko3c2dLyry
QGqBJjrnL8j66SAf3GQQB+0TdvyzVsH6zeqytdSslWrH8v5Gw75nqLL8j1m5aROvpFhJ8byovzbQ
7j0NQuiyAFpgz/OVQwCA66WhdE7pbIHWOLkf7P4hzBOQotFiXNpFLGyMKEppI638r4Zb00cpFnap
bsoHC/YK5HSlNKVs0kAvtlgU1+UcYiXU32OYVUcki37hatcTBnG1yhVlS2hTuQWdYf6ejntjsDSn
b0o/+plRqJDdF9nTfBfLEEMEwuBmMsd0/Z3VldIgsmM7f596fRKGLi7LBjD3VvgUDwQl9UEVzx78
2uQU0lQDefwXnkIErC8OpKIqadFGmvYmO0DfoZKC3bXvrKB282KYo0iinXghwJ4Q0IcRXiw40WVY
wOzXyj2GilAaHSgRHmldqFoX95Rdtz/3WUOFtlYi1moBCni+lZJzsR49BZghm9Ej/dPrR6JeVlTI
DrV2gKlb1eH5Ar/PY2RIqC1YBTvI4bEbfyDsjDzFQFyUGiDfGirMtwqElByytDsjU16UvFsy07+4
8KECKdkeoJCifkJzu92G6ClnO4MoyKl5x85hQxnes1MpdNBztdo6SIap9eJhcvFaP9sHVIBeHDBv
7+PrBoRrAxFXeetVzKUWMLF+IIFKu5svN2xLHixTeMa7syiBUqO+v7MbFmUjkXmPxQudKrW/DE48
jVu7HZky2BzqBXCRBHeAWqggIMnfmj4967sQBuOZm0UiEvwOjwXxR4ldPljDc8t8Yo4H5SjgdNZ/
E04yxur0uzR7DF7dmomkr4sf4nSL9jq3/OZa9dTljIwal4xyueM7pe7LQKB1aNDAvtGN1SGgTpk3
mLdTSNnxKpGCRDfDEYCGTSi20EisXq1ES0T2cBDWJax/KD9BWwUZSJQAVM2tdOwxp6u+k3l06w+q
xzqsT0e5HXOtqgtPu6L2eFueXquLvC0bHuGfX2i0aGmrUwioME76lZhe3hBwe2WRGNKq8X300qZM
E+tAiInhFL/cORWgEmXG9QST2BUyAvkBVF6wsURqbrPJVjbT4hhE4deqCfROxQsjfwh5acVxnEiu
5pOrE7iXQrep/05dDTl+I1N02ZpS577fJkIA6seD5gk8hkHDi3L/ODxkeBjEj5hrqKMNzFf/7NLg
8yb/ap+E3vGECBfzEJnq+lCW5bUPRl9eCsUFcPlHWlvD7uArZ0na4g7Xpcd41HQimUiIRorqUkMs
vrvwWX49j6MM9a4wHrjfFx4/nxq6hr5dOCP+DRbeNEI3L8dhbmoGbrHePCa8RI91S1+USDZ+1UT7
JempGRIxsztEliKxljsgt7jdHqWurRS2VOL2XGVw6nUSWw7/hEMUdF5/EnS2A7F587SWpBqgaoL+
Tca5Q3/1QlhpPZZXpaD2yhHLR1t5zh211sVXmLB7uIuVHNs/mu+oUkGY8pr35xLfRkpjpwCEvFUn
++CiWoi7RUmkKopTfl0RUyjKUV4KF0unmdhbLT4IyfgkVnicH1gCovojlc8Nu3oEejxFc0B6GhnI
nm7ZF+Tnw0WNjZ08f7GOOD05zcigd2cG5Uj4qledxIgNjjZunGSyg2DAuIgE6linSx90q9oXRaCZ
IYhfyB8wQnbY7sYfdzyvKuddCj3BO4Cs5o2xT7qL9oon9ycNDJ8Uwpv1ve1rpPupUKT0S4MkKp4i
1+oOGEHZY+2W78qGdQJY7Ghtn8kYlj348t257kUyxUx4m/w0JsONoLZZyP0u7YGamy6kGHHG1ADW
D128QkgeberL23k3YZ1gNXbxcIqFuVFPuZykVHbER28X5J2kX4zzIP9Bpm5ioJ5qIou7TK4VlOUE
EDSWkYWE9khXuUbsPJ8BTQPgLOG6PpRmpEjeL1QHSd4e0KPgc+gk0cqLYnp1bHntrn/+UiNn4Ukl
C/56oco99rkmE4lRGXlf1aYRcdv3RUbzWBiL/ugStn+mo2wjm+96nme1fK3Iyi+YwhL/WFUN0JZh
KvR8z9UkpbX65hVYWZZVeuSsRjCXcwD2ETlxxPL0X6U2JL7H5jQQ7eeygnk4HDjFZgl/zrellTtO
qOAMTJ/ssEnCOWTbTbG2muBPJeaXc3feNFkOvZ4Zdph/y5KvZV1/8jvFD2vX0X8ZtX/MjT/EwAt6
UeQtoNbi6Xu37SmHtA24LSTiPE/MSW/uUI0ueLV5B92AorYswG0d2KYIcXnkl6+981Pj9yAj0AGb
sw19mRDLw38oMKFmKE872FTyBUIXQPPF6Ghw5EhoyKn0nC560kWAFxrxr+xyvqw8Z7S6Kvn5Zzyp
pwXmDm/qSIogFS4JxLvtI04n9F6npdSEWycgZy+cxNwfJHdu2u4V/FYgYBqsx7zDjsNY29j8rS+I
tJQzcyWU636h0v8IkB06xeLwviL5WO53t3nBx+hJzv1UXFuTU9MHJxIZbAEPF/4otw4d5fMV57EE
YRkELL5efY/UmGSyLtWC5tqEFyvt4iF9vJZ/DcqXqYdZhhiiSEPR4wlCSQrAjus8VUJosMFcTMN8
/ft5u/2BZb7854ThboIXkzubppwimY31ZmJnIB6G6z2JkhRUFeF7hZNTxCpBKply0Mtqqed/Y1AQ
YTxMK3kWuIaYyGc557Zm5zozPLzF3F1byo12aqvBFrncKsvnKyPgg3E6CxmvXJhHz9dB7DIfvaJz
sCv5vELyjgz9ndelmbvtkrddjeYoY3BLl7G+iVDF8/0wQmhex+7H2hekg3EN/Ru9fmNx/3pka9G4
Yeu1yZzkPTqa7Q16Q94D2QCZu9x+5GfMJaJFLYzDBRecVUFJKtlg11KaSIQ84nq7UmKfjfDBQcCZ
IOZ+VHVUAVMe+fgeFo34UvhNc1zjYl/MP+SAfth9hGOABfKA/ffKfkKgU7GfyLUxKB3qoCOH4EI9
FjRQpSwJvAlXs7mbfeJpV3lOGaIPIbiSsbjDwRRM5+gwIRof0tR0swRPnDQCllrWli71CU18HhOz
G/4yQZbaPgi7bI9sT1OEMoYNvHprJ4cdMAQ8RCcMQhPdlkekJqv2CECgi2nQ6eqbYasjceS2t6sV
fTUnUgg7tvTbzmH7b4AKhNi+Aqg5nXFyMxZJqS6+I4rKNVVDlkuZ5+ZrGEWH0q7JYV+raHKZsqmh
qkn3sMikAunCuhb2PjMCKAQxe6/1SGeuRVnuFwwpCqbJfdYAOEBBaeQMPZw1mIwhnPHtSF/5r+N5
A7hMj43nIy880mdg/hUIQBQNAwjGzDSpVKaBQc6Gkn6qkVd0Qvse5Z0uOY02cHq9NyoVJdzWgXJK
1F1Cx0F8LcKzRTUyxRknq5W+HtsHFtAsIa4UznFqk6gc4I7x4OU0Pccnte8TNV/53tQ96WBCHaZ+
aebIckhgc9STe0MOESLDhnGvbDpOAj8I+Yixy0Wevl2zYe7oiCS+e2FuabtZ9uNuHA4KKk8JzY7U
DVdis8io4CJkohe1E+WOpKfYqA8PKnFI2GEadXVRUQkhqQbnYn0S63xX+5RwOUUYSGIGMICBrLt1
gkMI/z/Idrc+pOebjMIo0uStqEqUnScRhjsaY9n072fbj8RoOPi8dk0RJCyjXlv3SZeTgWEYIKOk
QEWbYRUQP+R+9a1FVbY8YYUvxV7JAwPCDbmMpXabgSaWRU1JBN1XvhP8Cxlq/W++gf+OO6Ev6FgT
BLnYbN3ooJAbSf84gZLzpw08Kr56K0Qx8GM/UJ+IRaylGYB5nMULgTQ5W7pP6NsrRaFxzKg+AfMK
2Z/gD+fSWPXzOJ07qZozKv+9voGjZ9t1ZWaQZu6qDkfr467CaXIITCPG/C92ckJIkXW08rOQzqdo
t/tRZQBXuQt2ph7irVo9ZUFh1Vy6+7UZQ+uG6J9vK8bwCo9Fi6ur+RbRVKyMvZdYwfxtKPpNRSPN
k9C99S/7D4z0jxQCVj0wIBii6JqJpstt14eri0saIEab38pEN7+UfNHl3o72nh+edWVU7h6Rr5iI
LIh9c4uLXGviqSGsvHBmhKTbo93EZSm1DcdO9f0+8bmMORGdX3LkBBLDTSdT9H8ezSrrD7Pcd3sQ
b+rUEeIou1TjeEwtwPiJXhpg7i2unoqjz6bGB7+uKJ+mu8NhbXjjE+fnLKF4oT6YZ0kitQbfbeZF
vZdRnANhtUSafAZn6LA2GKl1+Kmpi2SlFsGBwzuvs/danXmZEM1UUdleTrXm0LecBKV6sCpH7zP2
ulqiZoSVXQcW74yXes2e8v3GHF0r2M8DxFcBoN2ecsMDK4RRGH7XhLdhOenaljjHX7Ffj/8ONpSo
yqS+70NSdJDy/NMIQkJXjAauZJU4k2MdDjUkqcUCbuNljxDQWHoYMu9/hsaBAnBjZuwJZ9LGGbrH
1aJjiyBupTGyaiN6DytHL5BB/QGWbgtKCqlcd9bV/iX6+H9I9FsuSZ73nhlKPGeTbVNNQ/I5MVj8
HMGy7tw+wXrgCEmVPMMZaxE+xBFvl9bS3lQ5PkffbyFn0kfDvRrBV9XjgHFe4JJYn6jl3zoXKmjn
P6Rm8x9F5hIrKCcwzDBlzcLklFnGJVqB65LfbGrdnyMIp8yVySbjkEY4Qo0V1zq2VToqd9XeD4Ly
qnAQA/0Zj+oM3StqthMVN/du4lYUvfdJVJWbfOV9+lsPLegRUN6RnkKEdo06GbgMpyZIMIpjy2Ku
onZeOJ1zjOXK0oRiVriy4tCdhso+9ev3QiaTPHGhr2m6VF8oJrJ43aYK2ow9/rofQ0cVoH6PIsFV
AMH7WK+77U+hLagoJR7EYQt33M1q7zeUbqSrrb5mKV0faisGqtFLTuf5ndCnv25X4pCKNLYv0G0U
Z8dWfP8rqf3F406iH7Ume/ZpxP6E/s2SzzpNX516a72cbVp6b1CAKHFtPGg8vDXSs+ZdVaJ+sSdj
Kkbd+Xekri9eU4XYlqu3cSU10bB+2/rezm611sR4Z5QB0xrFJzwRscyPq7g9IsQYHkO/zjujyHG/
D+MFRrOxAbdzUGz6p8PfX4m3k7UrdhbCrZFdTe5sWzNZd3e1FSAiqoa1c6oRIHeNLWvPGm4O71jX
yA8irZ7NMqrK+uzzYyKSV949FCSe2lBOTnnbAIV+IkYnGQai0X1TsSaNz8yu84zZem6UlDYyfIcf
723i2t5F5oTZMpDCcpqcrjZa3eCzDHSYn6nsN0RscYXjArbQ2WdRvWNuMGDdGBCUWvWA2O7Sv7LN
YzJrbylPViUhhIo7aTBz+WtgPKzw7m0HHfQbHHf4ENoN1HEkH2fVJqDa4zKII97IqskB+BqCBo4T
D4v7d1EvXDPQKcx7o+MKrRY14LI6Dd+g4a9y2a2TU7YHGIlmjlU9JsG8XPdcWMDm2ozamIkyRfUZ
0FH+wI26peZ+VQyEolUUdqfoZjPMYtox4xaEvLu+pRUzCGroSjBrzV9eqfCkskdl4l4Lla17MmcJ
9XmEvZTQxBgPzCZidnkhrk2tqBX9F3i6ShDE2+CfqM5KWQC0uI1wSfzkeB1iHs8OPbjmIhxjsNGT
XKmB7QlyZb8RrZNoxskVWJZCOygP+qKOCUiNAghCJPxvX0kLlp7YZBFAJBCbU2ISWM8Nsn4c4M6p
rQ4Cj4UoVkfMTH5m8CHNsIAqKoCvWIs5oAjhI2iQuGDzG6Mjlt9x9YekrJGAA9psWr5Phgp5XFst
HjHXUzISyecfCwbuzWOLN6TMclmODJIJlDidi895LVU+eTj1WDFrMZVenz3mnzc9sJH+SFnFj2+d
3YP1VfXmt3AC0D/oOLECdD+zmq4e8t2oyYyyexiJD9V6CHFPSIukvR/2he1zPXnEKlSIVdyaYvrt
q20XlURuHq55Mxg+P/+7K0Wz3xUUtludA6EPyIH65WVZuj/AHVjN6w9D9xw07qaqLnRlsg529Lrz
h3dVoV+TdswqEf7Tg3/w+6tk66UcOmd2+fRuG1sX3crN7BDAqngP9Lek+Yq8auQKoI91tnYTbY5p
weJbPXfwMrQCPPFGs2MNovDsew9Ulc3Tvw3P/B/tXn4GAyBm2mxrHWIsYo6q+oUKobputCbGbSYc
JFhwWKHrPXAF4YrBUPzB/Xxl1YtCLxrwPKpShJMAyzj1NiVAJVniWD7cHA1uTB7SciGXScbcwABS
tzVBGxRVtrRFilasntEZ4qIsr4qL0eDenYKSxwYNHbz9SwfIKjEVc+AAQptxd/kJD+Vp+AExP7lb
Nif7HcxZDrJKoYU4BGwf4s9GfmlACaxDYidYeRNmkqywdwbcNHktqHQwWeG7Z069kLj3r02kAz44
Znv732j1MbgFdbrtr3dnppyB7v2rxR9FxU11V4PqFZVrDyhjc78oWdB2yDTjwUPfAbppRUBopwUN
VA1c0Tb7bT67I+DhBVQlzq8R+RPHEhHeV2gILREFW1GQhNrFHjRYo40/Fef1rc1A8U6440b8eKEJ
LXHtMErAE0WlO08B8ox5o6I/ieQc6GJKGXTnfGHz+wpsBejPjetAA0xjC/s4eTM9KmAz6BGomCE1
0h29uAfgovHBojI5wbJkcajefHKkEDuuV+wmoOfG3IPmdfmmW4JzRWrrmh6TvlERdc5RtiP8W+Ms
z/WYVzAesUyUGlXTKidK4oVUgPXEgQjjArNOaFN9OXVYmyNGK1PZB2nrUDm6T5UmnHmcEXcBPpM4
n7D01kCiMuFXErby59TvQvI4DuUYWyUWXw+6MqsLkW5DF7UVUqlqiEfPddvM9DnP/xrU7PXxShN9
mXa+ObcFM+yDjXYaqglMZTbylbrQ2zGEEnegyCzNE3mRirOOOlqhItMSpWMS56c0EEnUJmd8UyiY
3VTiFUA0bHonYHZpW/tcDfhK3TRQjaEU3+bEWr1oiRw17o1GXx8wA0uFbQ94f7CBa03MwtHfJoYO
A1glifJVapzTgKth9IbIwMB/WRiVU3pyorCiFhQ+BkOw7ghyqicDppUzN99oF/TM/TQkA/eWTE0X
qAaWAQZ/yk6R/es+CFjW962w67wP9lQgqHMyTLsWl5okSUhd8m/ScmqPyJkVOOKi65iSZLmcBVpA
ASJwUWG18ShnABfJi0F7rbKrcBj/jt7Fq6JtyoJgqNKsho9k6u0D7w3LyOQhCeo5fgdAXaLtJ/+O
qbgEC/+XlmDOfZudVvEeRg4J5WGG9B0GI/N7M7Ph170u+G39gXPGNCkt2w37XFricIWntb27UMpt
f/1e1UYicpjPc0PMt9p/Svu5aEqIBQx3IgzJVax5lrGtQnHSLH8/KRNO/MJEpUDR/W1wszRWh5cy
gSCqA6ik8vyWe3Em+GZnyzAo9GscybUQiHD9qn8fdp86d6fMaPWb1wrQSe7r1tU8f62t6fBgXjwX
nhabHT77PUjycwhE8t3lTsFTqkHEkL1ArOWMW2KYjy2OAueq0cvWAqDNrE3tY2nZmbS2AjNuIecO
iRGdY9hWNjJFx+irX6Uvkueys62zQMUZM0f/PgWz5nmnFE+G1i0UpPTxGwdSEFdMwoKhN94RELck
gPwAiK0UFq1nnBu39fXsSSHm5dZkcC16SsR/L2YCbn7iCavMhno/m2548HQcRT4G9Tk3YDA+u867
4NyuQjRuD+OiYompOuVqDLOiwsv94cG06SmwwAobegHDpeshDFr33SiJAXsK++LMyEKwuukpiRzk
qFZWX/WDgxwBuJwq6cMmONDR35H8Fh2QCJcIcPc51M7slU+8etdgrwL7N2vqoH9WtvUHTbP9Mrs2
kxqanb8j4pbmdBvy/T7+ryndOWJPpL76G3b4qGInDpyJ2eu7mtXwhZYWlrCIYdkvYWHyZKN1ozBq
LElNScv3TLULkmrusMcYHTLQKwxiRhhCbQ0seVgEADMdMnURL1GVYhANkYIJVful2474MYLtUDsN
aLEUDo197DL9Lz0rbkq6pSkbAmDFXNMYOQ47gncR1BIHid08+FVkCF+gVzhsr2eDgAuGlTtgrDNJ
Y5g0XBey6ISZuFywMvLY/p1sIuG7cKaOrRX80C5EEeKUJrEEz3ECXjDsC3UScPgZyCafAQrcGoU1
WSJUyGooALtkcEvlSKoB5n3m3jfDjgpiWM94hgx10exLFvntcos1AKro79Ri6pyaCRRbs9EL3Qpe
vyJ+5r3K4drEzrDi0iTEha8tm3n42qWNGK9io3yE1M9dbPM8q/v6I7M3cn+woK5jyqftNvdYV0b+
AhVm9i/Q7E8by+JwffC2K2/YbDS5gphYyyoCoCpwZpblmTahgjHBm2iF90Rv0KJv6M5NY/DcT2PT
KzKIsrq43HVtha6Gkmss9qxNkxUNFpq19srlUzL7n3iYzsB376X/LZqZWtfuIiziyrToj90N9eXu
9rKn1SuwSlNAyepv1VFxGFLtNPhmcFnI2MU/7DwmmuySTZJ95A4iEM/ExlDeofbc0ceuOIQYAQX6
79Fy46lSXJPmQsYDMYBOrmErTNiFZVRtPGXTYq45pE2VdZuGE3kqVocc9KLfgEsi8PcjjYW053Xy
1FMqDlRAtiSGeTq7DYAAIWqUu8CXBsmgzSMZlRNgcuClJ0c+YpZC5KWk0pyEPLRdn2ZUHBUAxiXu
DxYkINY4Eji/+qN75g1LLEJ7XD/I+14PL5oM0aCdBE5auIzV6/lAms7Sph12KgLaXSIf/Y9vKqb5
TreHWFgWLnKZKW7K41XuWYnPDxBCHPtIn7G57yVsUcpKcqggeXF4PkZY7wADYkvIK8JTcJ7iK6d8
QeD+wHh8z5XpWK2ZCy0lNBAcKipvwYUb0Ri7vabkC4C73BH1/B6+lELHflZL2A00hmGOzfDe+88V
2cNh7Diq5Hk6Xbm0Vc5YXMb3xQJSGSK2+KaJ3ZOZczawxnf/o5YRHWzA3KHXoHSRyfe2hEJHGLT9
qLOKScruh8q3oB4p/0R30rRVmMvKQ3gvXyaWlOR4uT3yBCXjmYSsHalq9pnuYDVDy33kkF1GNVXV
foVow0FQr9aTgLlge62yxdaKHva8/LRSacXzq0JUzEWrlvMcAtSLllf3a7xT1q5j4EnjHyJh6upV
cN3parHEVcQe2Rtf9PAvBtAZ34K0ZoFM7pB94HShuymzrZ+qWard1aeeOJKVr8zquEHwWxpPRnsK
/4FlS2SUxAAT3LVNqR/+tkTWZ0Sa/NMbHvbIPmCSQnJ89dzv7yye+Xa48hdTp+Z58/6+WDzDgmY6
baNa8HvFpDuBW7fhTlxxfosPqYMMKV0ghggoeTJ5cj1Csf6s/8iD9xpkcDxXqwflq5plgwQ8o0Ra
wMccYunRTF7un1/dHEC7aZEZrVS1wDHxIWomisZRsSI0byL55oRquJL79BT4FesUKxmrK6ngmxUN
w0FzvBkC4sOHbkQE87uIk9iixnyDWJW45Kk9e8bZFNRiUuBApAnsC1t6+S1JsQpDXl/MPbSgtxVW
bp/ba7fNJ+q3Bou4d6PdBpsyA4+Y2n1juH/T7WSiR7MDvDtjXyxd9Bw4mdNc0RiPAhzwPBLzaK5u
GaGUwFbD5Ha1eSzxEoVhcJaDI+X4XzSklCfpdpWMFSmNUtvVe7zEYhE8G3JGy7FTSf4NKRaHeADC
KNO3qLuGx/AM+v8vFf4ifNQb/nCyPeNBCTyGO9lnHBo1eu9HbAKE5cKz1bpjrwQaeM3U5Fpjjtop
9D9cB9QQT7hbkRUbRKCuQIF80U6khjJzL12legA2/OWAaskw+17VLfJ1irBSpK4iqfm2cvFAVYNT
yDy/0qXvDj78pEEx7d0X0OSx23bvlgv/MbapzAxCE13lNch575Fj/Pwm/mDUuAxgTsq1n0VY0yhf
eFtwMLWyUQtM5I21vv7dJx0Bl4WLxhIIh8TrFDj793+YPYyhwKhjLOq4dxWrR7NvmGMpo8Z5/zQ3
xl3hq6t/QdyQXrSWrZ0a6dY3JVKu7KlKGETaBwehYqOZLoCiA4smy4ln4k1O418/EoDonbYMDJGk
e9wJsef6Q49lwq2TnxcS34rMLKV1JrRHHuxDkI8sk5RwH0k+D1gzQdYPmEAEj+EtYD1j5V6bg+Aw
xhVw3JF2211yHyuXW0WzBRJK4oHcLceKyh5hikoRYaKxMNedMPaLUTQY+VHgYClPkSflmhjuQwK4
nghvgCxQac/BooaIQ1K1PwXKMeLVFnS840oKLtYZGsZDjti9X/sK4Nf3ll/Eq1LJZJhJlNz8wxeW
EaCecDEw6Ms9VBUHNO8vnPyThHqF/1GxDnlE0dLLON1mBmNgJy579BxjuG4dy3mipNNlAm0yysKj
SUHuC5mj4x3QOitoqdXOHGEaoVCRr0w05YCFMymO+2j/Ga1ZBtbYQF18H64fbiBXoN9hXg9XEJEF
ljwavETe0FtC4SnYagiYQuOtxzDZ1pxubKAlFkCsIIteb5QkgwDy1KYZA+yJDZO7D0wxv2ez+oZx
DFy4wHFE/06iPMOeTg1cTpPbQISnSxt/hZqqqIGA279WRt1bpAS1CQM9PLic493FWuAv/4YBHtK6
tUvTP1nAuvmdKncSvUQry0BQhaJriVl0A5xhOe/l+eqgjtomaYqU2MCbu4SB0u2/zA5UK/H9RH+e
ZiTUpe3Ra6sMuV0BnIABX7aQS3txLZzBl5dVm96fbiLft7RammI2m29cDKqsxBa81ITO6/OURCD/
+FDx3wrJDijjI9bgCWUaZd7gyP4l1MBnKe6xgV3J2EIlHCg13GoNtC4k08ddLZ9EAqje0jJ2TgrZ
Pl+L+gx/FBUN26rfXNFOlCGMXO0X9+jsQdkflNWQIM5xgNvN9LOkuXh0kTqJLOh21cwy4wb45BRM
X9XF7/Uk+I/B1bwYNGJT+F4VhESjMbhEHnMvsTVhTRyZFNzLfEdfuR+QaVh+xjZP5ySXWssfirYm
ZQte7soEwqPtjhhD/UmnFGq6AClPi7g4ENzU7WxSzcf7HY1AdgQnrdGBzFjantV9wGVOrUP96/H6
sKg6ESPEuDovfKxNKqDtUBzz9eRr3SH46HhIS56wV+76yLocvkwQ1yRbFdHoI4jz3Dd2BmgdBDIR
LBTKkxSUKrmPdi+ioR1F603piR2KCsmWipB9q7MPa1HI2jx4jSpBQeLnoub0HWr8uQT3bfawoNgk
1h4/LYpXKUeTgpzRki/96wD5hOBDB4fwTVzGJbvRLBumcZxzIttPMVw6PVVZ/+hCplslxcF7c1+J
bYPaMFAMIXxOFAHgOReYvKd5IymHQ6D6iviAi3vUoqrs9NAhNe6EIdaFhEvV29mfCmVi1JNwugWl
DpPm7wJyzUaLHpQO0YJd2/Lffeu70ala6Cpc1jWZTnH9HudlSWVZNgc+I5P8PNfTm6k6qkufkRcl
p6bfN0QZRDlm+pj1fd3gUnwbbp7gZxQQBwG2hmdlC3p2CEsNrsadndqLMb/JDk7qLRqgtrhyZMhc
8jBp/8bnBsNF5aoSS0CCHnoV6XVNUUw3Vjad58z1F9DMPJ/ffMFOK5a/SiWtkzttSu5nt4xaD3VB
UxGWfxum+PLgjHiQtkAVUaZWRa11oBXILyIvy870Wxo3Zd/LXl5NqBrO/prwNQulvlqxciLQiyca
a1j9mUreUjyEp89frGbxPbGUcNtuj04hhNIFVKg+Ku1XcBG2CKKs5FEDGjJsPurAWv7mZRkDulPX
vXe+w6/I8tiSQLQedX10wzTEikm9r8JfBiFp8SXehpwj/Xmje9+pkV2blk9kpHIcpSpVvCBusXhE
WtzmJNUab8QvRGPkYiekP3HW2jrDtHP0KdLnXCCfznT8rJ29iZW0srJLdTBcJDmddNJjD1fhjYOU
GBV7gQc1bc9CYgD7EHpKmi/n7+baDLRhZgPNsj7C69TLRUbj70khRIUYarT9rLQeRceUd4ZqiWXu
g+wFVrAVRe4a1tG9vOOvzVRIF4i1oI5MKBIeumU9FTT2W9RjhbyQAI/KToS0S6138X1+TYbBNxOo
7sCJ76l2gtCiQ03MemtEYLHseyfNFuh/2TGUXxfWCc913AngsB26pXqZlLVden8liNEsM7Mj56pV
lC26JP6SH/jxiZAY5nHjlAytie6KrPodJLDn8tvryGQOtkYgZRcj31bZorL1m80VR/W95SNbnkSn
2hb2QSGf3hMvobJ0aZ0kh9sgJEdKYHuyV9fFThdf2VQYaXm20Spmbh+PnyVGRZcnrS4voCsKwa7v
e/Zj/o+Y6Ghv+27/o8L0MA5+gr6RwjLHEsthhGo9ONWRFU5TPadz9eSDLxwisT1nR+hx5LURk4UG
FOQKXXl6/7MWqQX4jBPTvwBlmPTZZi6CIKpZ2Zd3vleyAKkmhdp39M0+cKjeXxyUMtGXbRkCPx5C
pXRqOOWhPRwbbP/l6p/7WojmANuZvqGkkXcHXbnXMvH7L34s0Np6caE82HxQmoUfFHAHTSp9dvFH
MiG1jU5J4sacDtF3idO9aRO38P+ktJjfuyu5WmPFTwG7ZrOIyst9gp9kBL7j2s9yiBEWsILdMTog
QZuWcN2dpfgfY5NjZJhBbaPArrDxsbKUUjg1k1zyMKnpeHox1AkMIi4P5UHVe+0iorum2+sBvkhh
F5nowm6LB6kA9fp4fr3UTZ5eXNwB6k5ulyW07vsQriAYZVvuQLylphwNwtvaAwaWXbXXv9i/Aig/
QB/CZK+xsGzszP8mlqvNNfiwF2Dl9LBvrHR2dRca++SrmeIhYHCjNbjVk2ui1Kdd8Dk7V2MmAIhi
3wMnhKRZ+1u8u7mTswG06of/XnNoyMPAkjfJRWvgaut5N1CGdBvgPqKmMug+EZz5en6zgorPBvXE
cU1/MlN0AfO/jqwIj3d5LltOOgKLrhqhHMN/9f+chV1YS1TFsIRMio4eInZcesR+lBsXlnlw0iOD
v9XhN8uvHm4GoOY8YmVq3na6TYNL/gy8qDHdoc9sGQ9udmT7Ai6LrQ3/CSuqIhX7mwZg+D+LAHE4
8/oaf3gECcwFwAQSsW5wwSIkXr+MVNNACfVBzC5sN0FKAAHq1JXW6sjXPqsLUvc/7NYe6K7oOkcs
RH2IvbrU9LW689l5bL1G9KFLipJn0EZkWVc0z+hO9rLAoRl50dVoume/4pxS/14ncn4mj7Nf/Udi
ditdvMIVQidEIv5IeqUs0IsXJLouDgL/zJUfIY8EqttqZNomjgE7L7UyjK3iDXH2fOwZmp7gb9aO
HdoqdfmqlP2MF3YN8++Wx46yT6GpdLrAsUwST6uU8SwTdEx6ME6nHzhFbTdPdF8IFOdSZsIzJSWn
VsQC3xvt4cOTwJU6Eb+l31hdcOzSpTiAa4GgeFjamR+5Dn+yniWRk5lNMZqB/D5T/FmhBD05oYA0
FMUi03Za7tuLh3kc1S47pUTTENiYtH/vVeWCZQDvUsJAPlgZM1RkKfApOI/Ho521nks4X+hAENWR
zI6ng0PI9fvqpQ4sGDMLl08uBifUFO1AioMPWS/S6bPsmpsKJvcAMSk3+drvAOPoRVdBPxtwe6lS
G79VW6I/gPJcmOiHqnZOuS4bXDGi3Led/2iUVDkt7JVkjsZ3wFV6FZ4N7Y/6quBu5MyDNkNTqbQw
w7T+jSt5luAWYNsjqy2O7cgycDAPGb4u1dOcOumT6WdUZQmh2wdI19SwGPUigFe0W7TvVTfxcgDd
jY718f1/BxCTOrT4ijXEUjmvMzYq6+OUnhyNVTk/HK1WgXQIK7z1IPg9z+TBz9wcouQc2i5IzzXA
6V6VS4OTGDXav1UPn/y7IVtGxXuaCi8VEUspcMaPYFbnr+A/M0wIVhFjmJ4koqDZqemRvN6Nsjcb
+AgUEfB8rBv/V9tVk1xURwoUvTZqkbN+ZHu0hQdIjTj1OwTuYvBYVxXA9DdDS8Cuz/ttzagLmp0d
a8rpeIVO8ALtkP+1eTCCpySXA/ftQtdZNtoyM18n0JasF3SyWpquomssrPFfDja7gHmFqUJazaxr
cgt49JTJyumTEdek5MEEO2nWMt7ep8cs4vBq5pzr12E9yJXRUoGnx+XczZAh5AmKP1ydevqZWLjj
lc30CiYrveul3/MeN9cHi7pQfKRu7hlsrsOR5iQbx1lUJFvxkzOgiukFxwWUP141qFBJf/u03tBK
ErIPh/joLz/w22aGNDQ8F9HWxEmEfoEAhG7AcaiMG6e9h8kwa4ApTKJ9KqiHNp9RliFypEsTKWD1
5WX4KUrYOZwu42A3YBVSvce5eoJ0tEbtBo9P9s0L6DcVyvrfGUwmPuMooWUYgKlpS9qvZzDTGUGc
rjJ8AlIb9/qE2g4kBBak9F8NUq2C/knM2I6JtGVlCNPUGpeD0TgIwOd2yCUn1y3FGvkfU0zOjvwo
euShdfZteTJM6rx87WHNkdrDuNxH45PP7b5wN+jnZZGV2KNy2XFDroS4UucrPByjzgTgvdsUHdn8
adb4mUwekO0LvaVE0RElc1ekJE2fSxxuQ9ulKyuazUd+FZ9WOvl2hWCi80jH4keu0C/u4sbw6POW
9NGIB5xh2/v+B5ODahBdgz09ttcQ0uTFGFEqlWZFQPy9gqD+31NEl4YoRQnxt83Bjt5nMehFMyXo
XwjWptQOcSRY8G6QGriGl9ZJiYUtCD8LwRamSheV/ZfGFuu+mDYiNINlB6qFnmvybKc0F3MLfTty
e0wn1q2DOPxYHhVvRQXyTw/GZMUu/OrlXP2meN+TF+hFeqxA2wOClb4p5khX5E7mlcvOkqFt1D07
YnLG7DB97ucQIwqOqrATgr+bb3KTE41eKxy3w1IwSVWRVYAZTLsmI24BcDiMN8MolPYaObjxXOKo
lEFO/fH04uYzkbQwD91YMm71N6YwTZPkocZZNkx93K4gDbrpI0QevBqLz8L4xWmLgr4TuI7lBsjs
WsME64maRHIeyh3ZxXx/MLVPQWoEXo03B4Mm7kcYGDNqTni4hoqwo8IcPTp9QU1Ar17w56NkcWS4
COr3obTZBcNl67PArmIzA7k9k4WZGqm/R8Z2829qNBozN4HThuC5s58ylI4bMcmV4f6vTfTB6GYR
SnwY8T5W1CADhhFKw/+ct7pwauOcu98/GwC4vPuNMPeWO9Gq5a16R++CPYAH9U7nUuInrn1SmoG+
5kf9P8A9UY3ww3Kje3nUgq9nJeuIFQKmNRqk8CWfROqRMxzliuNCmTTadPQxVaXrIdudpaM4Uo43
j2l8egRgu2ghtuGy4LxsoJgoNkgG1QTNuTZHKciIBsQJs4/BSb2pGt+Pyy9Qo2o36yRkioDo2q3n
3NWxo1ky0jbx1xkcZnDT7p5joSN+wy6fmiznifg6LXrK5aJDznWbRkByKD84OyvzgHPdR9Nu0++h
NhmEeoealGgTojh2WVb6nNKZR3naG9tep6X9D7Ha7Y4Ns86zo3WrvBeJ4LfDGkc0jIL6Wcge6LhM
67DCnPX780q7vmWNiGRfcqmtTECK8ZpFPb2xY5RsrQ9VXbNhgJbvADLWHfh0K7HqGHfYD1hj8CXR
CVPNxq9U7Ul/oRuxWZOPWBHgV3QCwvgQ7ukUc2i4VjBRl2JcV/2RMjbI4AkUwQh9mMWj2gZNxm2g
oEXnQXzXFLqaY0DnQd9IOahImVCd18/6ax/mmwbgXCgwqoOIjJF2kTfoHStpksYUsVp7cnu9XHq1
NkyyLeBTRRFtxKns7i/bJB3Nd296hgOFaGX0vpNXK+3wlxmPxCcoDJgCoBexw9e3kG6qoBvWxIJE
n5MwRph68U4qmfGXC8HlK4AZllbMoAMSgsgKBOpIrs7hlbLS37FTX0S7tJpJm9/B6xIjfkMj+eJW
8B6qRVsvzZyOfli4Mjk2N8ym9QuotwvnDVXdmBiJzGT76/AHy3NsSnOQ61jcfIzU39Qy65uMyGCm
ZA2PJ3/gouhe1OqfuK26ZcCxKU080lTA6ryCGjVqHofS1jjXBf9odq0ldGpzhPDf+RE50baRfxuC
EPzhCtk+GP+ArHBlLT3aqvZvlZwZoiFAsE/6sdg0zzm8phZtqlWc4+psR+ojI6Hgun0j5UQVn9xT
r1ZZ27cRi4HAZhgT3A5MzqpF1vVP7JBCKrrZHd5PpDZbbsn203ms3mro8PJ8PE5+/TNyHud1dkKH
qDgqyRc7P1MOKyHaf4kk/Mx06VFAK8WQURC7E5OpyjrJLyb93eSjNZ+Ov3hqnEyO7fL5AmrijNXE
rAKWi4lq24HYt8nD2tmTbH7eMS1bKmqQb4hbaDKck85g2wU30QCAKCpBdxVS6caWPmN9WqeGDwAl
bxWW6e+TNkm/FO5JZCZhFINFrxrKZ3q9jB0VWDaV5HQnCf4AW49QyyJtizLkz/lU7+MGu8PDhXrZ
mIjo+egoEYPLotFPDG8ll/ZF2q70vg23KKRXr3XBGkmapX/gvcOVZ1H1zF6ik1YZ28ZBT3dljdtJ
dLHVtAvjSAVsY+tR+lU36kfvSEjqEwYcwNoZq3KKejxPGBKj/r5411mZCUTlk9VJnOjcHLEYe9NR
ZV5KKe6Iyb5JmNcZYMvsORfiAyUtWRN0PRF5v0UXBSuoPdN+E+dJi4faG7klmzkcFq/2DHAyTA8d
XjLaLrbjTSDMDJYH4hfzkjhCWdob/M7FOGzvaW0u4w1RpFysh4KHkzs4L/SlIIDCnA2pnH5AjJbB
/GLh//ijuVFfxhtVcXT7f9Qa5y/CrdoJG6prNf1bNprwQMxVn080HAV9bQ7xrrzi0JSTvjcLVgMQ
cjyR/bw6FFmTTpZ7TPcN/KEMnu+W12hqHDFUb05XSWRU+bZTEuWS4xTlPzSR1g58JuzdKfuzviOg
kM108ACC8vRQN7eiLzQ+2CdbC5LxMpNf5Vq8J5BefEjipvDBgnCHeME+V92EBpsuYHnEta1w7ftC
YACpzlNTRHVNz51S79ZHQ8+yy89sN/fzIoEmkDsE1VSPHpDC+Ii5C7kDCdnk3E7mN4fwy232fOeW
LLd7IKs948MEf14W8AJYVuLP+MsbhyAL/xT6JYWdqT+t9WYAvu4sc9rP4znw/oYH3kgXvcI+PSlr
YYjRbLa3VRpNNWbjJqyCu/DOgc0cHa5qbk+x7+cdt3PdXMNfny+N3rKbCZ1LfZ2f8TI0AqeRVfT1
q4x49c2F+4/Og+r9RBRWkFky+sLUk3yjE2Xbq5VvEoWnFGjPjup4B5WCbp8mgU5RxOp3h7KJPckA
fUOmjLGb/l6/0amh92FQJaUgjwvNvMsVkkWl7G7dKgp86Xu/bQOvC73KRA2MVeQwpMP63aahkK+o
DCHr+ZjKDm3EWnkgZIBWSVGRvgI7Nca3zy2b9uswChJFtT8eny6Dr3rgYEAD9bulbftgGlWtLGEw
5ftbH/jOezV4Q4idlcsWvbQVcrh3QvxcyfOWiRoLRVyY7oswtRXXJS1ApSudyfyNsT9YJ3nteSSL
DRLYMd7PUK7rWXi/QgeH7vcJdvpZKWBVXQq333lZsIWuZXUIXe+CqqDs2qQ3FwLCBMKarml8u9Ir
5hOIIlDDQF8n1qy5h8gb/NRGUQ7pwVFV3i5OV9X3eI+aLVVpRA8O5/lKN1p4QTka+Y4X5S2lK222
T1Sq9tSL7rnh/e3AqfHjn23cdQA8d3rLDPmgyQ/mq+YI/VeDfT8Tnvp3yXXBKK1ZtvZVyLgrHCoc
vQ/c+mQFu2WDhCwaUsX5yUa1vVX1XYv0W0o6vyUBmg4oCF98JUEujzT+mWbHKeKH7XIOXCkEs2B4
4gPxIseSsYAxSZFSDdePP3BzvbUWwXC0F+3dAc0yQba2nkxJTzq25ldITPVaMr8eX4BFYIc0KMZD
NH38kaNIXK6dm7UOF/un03qxAoBGD3qezrzvj5kcuyrwrxUVSnitMj69/Y9oE+lFkIRUb4eD8mT+
BOMwVBx3IJR5khK3fRtaKBSKiEG+9DUfGTSoiImhSXYrVh7X52Hq6W6hvGSsf3QksSY0KfICu0Ts
9ZBKt8PxPu1OyIRbvvo98sliOl4WHOzmPIolTQqw+z4jxJ9Mykd7wapgNo4iGYQ3I0wdo4HTIHGb
SsE7JJIy9jXBu1WbthkWSSQjhK4eGOgIkRUsy7PMdkJtuJ7zDizQdowVImrA5GV19kfFdiFQZy84
BssQzUgnhiw2PZuT5aeIv6m9WsAGCL0peWQ1OcAWJ3+kvDH9zOhm09Y2s33ewe//lXG7zBdthfof
Zp4Mmo1pDVmsHnJqCU4UlRQtb8/b6BfpnM6/GEJHg/pqNFnwHBA+zuOYTltl6nPQuqLDgjXSiqkX
vE9OYfPMeUKf5ycaNzPtZs+uEVl6HGERVt9KXosHf35Y2bTzvLJzD4OwTf8kBOPa/YhvldP6JCUc
e3rOcXAvk/h4D0U2Hq38T0kMko8Rh/XwvspoHk0khX7yKyiSXE2avDGKmUKuj+18UGq/iZguKbk5
9yDJFNdVyFWIWanlKWDTtya1en0ziXihMd2Zv4BBUDbT45LZT8eevjlNSBofY0VM0IddByZCqKUe
avIPQob2+OnapdL8hTjZ0KyD5VspbuuL27MFeRGID6RbCO/S8FUXxkwdWOBYir4aDVm0ktU1yfvR
Zbozn+tjqUt2/tw7OiYoNgFEZsPrtq4YPsq6Z6P/ngSIVkefN8XXVyPaE2kUFJ3ubQJYQlJygmyv
YlDTtQvvejQWriRtPcZ9K0eemK56yQhPfApIlMP7EJXwQrTK7LCqp0Qh+Wf4E6jqnik+AL0e/0Lr
47i01Dk8bQ/g+XW7crAOQk+v8+zaoF4tEhUZXxsoEfe72U5vmjiPEoX85Mh2j5duUSG1JA1y9OSN
M7LEMaFd4mw2X89iXQsl1SbFCAPFQdXOoD4X/rnowEYjcE4iPpMBYnDDIyMdAyRW2Pvr22SIUhq3
nTDVsb2jLuoVW96WvZxgBB8oyL+UheM8pyJZvF6UX5o7TTVZ2mBNCqZLnhBttDrllKMSj6PDGWm/
75wJZx6ZBndjrab+pgemRphR5fkjW3Yc9x6sMYcW1zLzL53So/JT1pqqpb3k5sGKZNn7eNPM1RYr
8HiPZcB2LWio/6ykwBR8zhkBY6gt1qwlGfjEKACyD+9ErsPrS+oe2E11rwwAmlltNP2KpeGspCsN
N+00039ee9dXjKzwgWO3997EkcEmRGzFlmiovWG/5B/pgW6AOJ7Xheyle/IydeotI1SX58GirX5K
Etx2A6aorwE3NqWgK3VZtFaUbme2ansoOvSModNrmJiBfsQfCykOlpwOjfvY0e62Vu7PNRl+apYH
TFX7atqLSkMr2rIDlRwoP+4SjaKVD0F6KWxIcSK1PdPk/BDlSsuTDH2PRiyoY+VxeGLjppjRVZGV
s0eZurTam0QIoEvp0RS+rKp1uE/E8+BHVFiy9oqzxNCvyz2Bkrr2qAwdwCfj21LHbdKai4V/qlbV
UgpNr+a+IlYmQb0bDs5AYuEWzGAPNtlugcnbj+/ryQ+Rmw+lBeVxKsJpr7cn2cjbaZ9eYQIYI8G+
8GIv0604Rv9OqccMs4MIFNw+bmPFh11m8OhUjT1OmWQX8qEqpmtQOKAkI2zNP1CsV3I42tv5ivxN
YF8uTifu/jCcBS0Mq8HZZEW48rH1JidbfkMZtrOTXWZ7vIqajenuXGQp/nR3KbR4bR7Svadqn0GZ
aQ2B50LKS1udY1FjrA8RjwP8OPOPIpwZ8YgT87aPvbhV3wl6AEaZA+Td0EtPueZbyDPAjOQW7tZF
i2nDEXLzWIB9jzlyk5SLzIryUC7Y7tyNgwSLAAmEjMwm6G5PkLXjSvDoA9Re703gwIFSmVFnapp0
/U0epRbQ+6i8XyAOUBAwl+0FvQYtg7lOvQU7dAvpFSsYCSB2NEnWyrrck/MZR5o48hFIrzpDGb2F
pesyQBQLzhuaJHid7XHbCcSldrsGBGHn5QO6z+xGKDr90KA+IccuE7YvqO1Br+v2W+QPpl1Z3ZBg
JF+RH1oFdE1MBdTeAfp7hVY5vth5csVX5orwxOdKrlfn/vZEStNmPoVqKs0X6z5ZmY0UON9wsMW1
ybjzsOusmWaW8kuoS87Ps6/2ZmCO2/sSlVDPX8MsYd4gFMR/WXH7P1i7O67xulfBwLNwSugLc3SR
HjQZvxQ5MTNorzRtTgrGpfE3YHIOEJRQZX3lqJVrzRgPUfx/IbeETX2NON70bjkwdZIrfB3SpnxS
vjChly+1UL1D5a0W8iVkXVTA9p3FNeUKmManIyilEeQfD39iVskVUtl2Y230U/+nYkGEdKizRbJz
cwmxY0xvlaDZ4/pejzYieY7mNE00CZo5DRHh+mwLdza4nQrqbKDcd/5jjCejsOFrXe3ShcVosaaT
WbacA1hWIGiGhn6R9nRm9mv+xVKJAAX9UUR3uEUjvMv5TRcOyehrUML/ew+zqcDVoDOcEu1vypO1
hEouo1SQPaswMAc6tGZbzB8rzhZkearLjUKSfedXOKZUYTxokN4s+2tW2X+VteWSXP676ZgAbb8n
4xZLu+dujeegE/Ve+NJjLMi8HF1M7nUYmdfo+J3ZvDaiSoept75CAhkttDUtH623upTHcD+0XWPP
cyWICC20djixyGRjCeFCoxfk7DXij15k60MFlE0Es+gfqcN+wz10BjmrbZxF+HStrqUGv+YVQ4Pe
ZMXkHzsScq2mdHvoTj4Z2sjKbRnj8RfivYVCgUyttjooOhgyK+d+jNYdJXPBl8QsRQKD/g0rWs06
t2J2QzPiDqCFIf6X4TL+dyYZyktlZGVZ1cWVamz9UOh2madsV+uf3MbyV+Lcku4+HgLawbPkLcZN
lcNgG7GZD1H3tlvkIM6j43+3oob0YzwyVE6Bw/6hvx6RR39QPLqygd1e6U2h6TTkPM14XGuQBYoT
MYOuLTN47L87zqWTca8UVUFLKEtwn9lPTaUxBqqjn2PIuYvg2jd0E4sgnzNULdcoBYN//C1syjic
kawS4+IcCHeCGyjvFDZDAL1NCOnjDMUY197k0h2i3NCbnuA4DUY2H9Pe61+bAmvrm4SAmVw7ue3f
IleLbsbF1NFD6lGdi5iXRQHopTBGfy1dG0rBNgWmZH4fFN8sXXwg5GA/iYAqnNLx0I6XnovRzEvD
63KMZ7BHkv0xez/S/tXiG/WRP6qFxjMIzPsVRfe/GUIXZnktF3EXijgVRO6jjRR4y0o58kMnmIJ5
m85pd5Pyjdn29RVhKLvUZfD4Ot0EmcNsZfjcbcdRYtlZvP2Vk7ko2Zym0ehQPDUfMBUqsrdWc9SZ
TpGxL5i809rGNcz9krjKuVeDZJEq0+GMsatOkrtfzHkrvL9ZlNJZ+561i0uP8tKeUjBaQswAPhul
wrvECC5UR982ptpLOw3IjV53n2ocB8+u3EuzWlBgrMZBQLgWWLeGwVx+J1E8vrsrLG2FBpP7Hrqn
o4r9bemIfpKgmO3c0+xEBHcuYMagpq5iOQ6ZuiFVKuThlxtMVjGLfRqHz+amPHkGe/y/RQggBZOW
njxvxM9uSzWhdeSPXoqmJGllUrbYPDvTOhHVON0UfXiBlKchucG5qjks6xCpMzgAZfpB3dSdtvH/
jNK+p7y8Z6P6ETC8Vjnq9VY/OsStaqjfi2bdAW+1AkJYSM7+YOOn7j38PpSbZ0eArY9O61ElZZW3
3QJGU53HtCK+tVpY5Kc5l6a6boo6WqBWfdU4QeRJyDzKOnZfq3FBaBtsiqj+zCM7RskWhejQJPdf
6/S7p9wQNhX79Be8bNJwwuyalTx/gl6I8R+QuDxvkb6lDurYWaEnKq24Tzsy0L4Li/W/jmICFgkb
+ZxYrPsr4yBoBqTB1A/WaVNR1jyouI4QZSWzrrqVxzzqyop2+hTHnUOO4F58INp9sDOZowyU0/hZ
GoCiOd54010qOIAh8Y+VlwGhME5IRNqDHXEXdYcfYRoqELQ89rwKg/qKwb8XMFJ86qSvzcAZCsPS
aK2WwK1YvE/kcy4ftEzKBm2yl+5ZjGEetKBuJAYJke+QNLTVCr8/TnLt1RIN/fsHxO3WkY/VAwUq
5e8BgWKDjB617vA0etaMWWWweEizmbNEFbeRhuT+dX1XBtQXHTekARGQ8Upg4ySHXw7VoXBjleS9
0/cdK3Cr75GnYW3FFanKmncWlgsn0Rx1tpYPaXwjcH0LtD6LXOKzOAop1jGqruKtaZA7FIZplLPj
tNIJxFF5zbR1as+/CGzVAAZ+Sf85f7KqnvwiIjk7dfn9k2ZMUqjjthgVb5Xe+Q7NA+sjxDx9GlMV
QtdBbW/8E/V+n2kPzPgnexBRl1swHn+NxGpc23MZOAU2f9F+u8/+ueVZ7olJZz9kO1ZEG1QnIrfw
pCutOMXdutmweKN8HWtjp0o23kpy67QLcpIkKx54XI15OT/cMmdK9VQW7m1kU9S7le0tI8C/0Vhz
1LeZGKKrM37w2NFClBysWtiIqzeS/2udpRlpMJ5DvF+iO8rzU0FgNH+UV6UExnxHxvJ4y21bIERv
Wpj4vSjM1JbcZPK86H/Hlpbtdjp9gh54/lYmb05CHoc0TZCSrDS+X8m9ISnCjl19j60dWRrqKML6
gUQipMDZRB+KrF9LFk1JLHfVTyJdVj4Wmtd73qwn1hlpxGQZx6fnja5BRdq/yFXWhDuOS3YkSqhm
Ql/dN8vVzxa2Yz2sZc6GhhrO/u0CyRhyftM423UbtY10fjKrSo3Ku8xf2yD1qIdhha+QNdhHlwvO
DFiXeuAdS8rv5YXPh7bQYG5oKuq8NaaCD2QhQOX+TcEjq+b3+866TRMHtjW9xtTmY9ZZMCuN9nxn
MtoFyD4szmpylbCtpqxKMiNqgvibb44GSzuW4uza09WmZGXDRctis6ezaG7JTI+J2r3YwdHakWw4
Vi846u/S6Tq4C4buUeaFQvm7qWpUNPj6MwdMcSZyCaxrmRw+ioqx0cZTUJVLmcaIoi1+pCE80rio
wX3lCz7zvigou2nTasUI70425d8WC1NCRcKi2c9QN/UMxoNTD63wBE1LemyfEZxphweFeLDe3oq9
y+4z6kMD37rl7TLaz88PMepRhP68dXLiuq7lmxEte8+aO+WnQksWYaB/fD7TER///BaLK8+HVIHt
kPNNt00o77vsnbs+Tw4O886Q+KrsP4Q7vlIBxgwHxXMdTq7LBdZP4YMmsYf66CtCWsfdfnjnQE/8
1ZODrinIkU9mwKYEJeOTM8dLozWM053Ea/90ewnDj6601aExI/Xhr475luuH46+X4mK0o22iRxm9
ZBPcPznOgI6TF53tTwAeMKJ3g3QPwNhbsFhb+Zxv87TndV6HGutHAaeGarF90Ce91KCSZEfiDNkF
JOpaChJFhIhuMGFEZp8MBfLs0+iniOmZ4NPa1qeIyKPQdybTy/ofNYrE04tOHZ/fVa2ZFKmi+RnF
U27NFZc8+uivpsjtLAqaZk84OPXRTHN3LhjRHTF3nwBGvq9T9nOcRuPC5frfPHwmLrNs1NA+lSLy
hu7Czraek0604SXybbpXJ1hFeso2XfM8fCFhEWjzhR8yT7FwMLPVLZ51ageGc+9o7WKf4uXVItea
MdEhXIxkPUdiTZHWJNgzkpPOS+nEH/R3cecTkug87fPoDYWEyMpqGXlwMNmKAbOuBod92K5QzqW6
72P+n79F1ZPI/86CfbNMRn0Lotx5jxy1yo7OEZD9tzU0LaE/Atif3NgVs/tDiaWg8iwWcArh4YK1
R8/c+D9D9qKOs4fFnC6s0BUyeubzxvlTvlMBfxDJ3k6mtqHWuIbXIRhNSAbu5j/CC8STIw9vJ82w
BrxzoROWDxFDWLJbZYzBjUyCkdmb7hhX1Y8qn7y1A4fOa7I2Og65OI3d0mzi5WBjy8lfhbqm/Kpx
ePEPJInaF+aGYOcrHaIhNYauRL6NaA4fm8OH8PgKI3K1hzwGNpDTsj6ONXSvrHmkl4k/DoOWwdm1
YGJRtIgq4JeY5RKMwtbtr0AC+EBI5erAlgs8n8d4+vk1MeK59yHclWBJ9U1feLDtlY1ywoL79n18
0gd7uOjdogFPBPreFq9DT0bNzz7XQJFFJsbNHY6HWR4CRspY3gmg9XKkXJEkB2DwEUIHqrTXU/lZ
/SWy4XhsakTS2SJ2djileBmysdinPewDPUzUY9lQ267dqPuX4WieL6qN4StSaGlSNotYq1S7pSeY
XPjkkSa/blzCig5Y10B6M4HH2vQU/fXoEpHHCmiMCOBWSy+0KbRUZlRJBr4YD5eI/SMQD6uaupJP
LKPTzUd7KUPeS0zi2FGs/wCHIBL2DF5Vn7gmT/yM52Eim4bxRn5lY6EwQ7AgFK5TrdAqRuGr6SZU
E63WErxglDfyF6pinrsUlijyMXCoGDE4SUx/PjL8TgNZ9fmmQ/wV9qqLCdr0j+oA/42Xsp+Trkw8
iRyoRgcqvKwdc3x8L8fRp/W/mV/WBJTu3ogdhLJPTGpgz1k3BdYmiuaw+hqF+3cURmkXvf7n6pc+
gq0410FAmjJ1u3PLnkOcXWC6KUu4Wkhafca6k7PwHcDP5GB18Qfo7nC2cAjU/DVQLSMvLe+pgKaW
XC/7IGZQSz+Io4sNgYxyAXF+urx4bZrjLpSpLQ8+6z57f8GDP3/EzBvybYrgP82UqI+q5KW/uU1E
IMizloQATLFik13yMazcl7l5scxOfJqqhIPu0RgPC4lBMeHdkSH+FriHHKzwzFwlMCjnzqEzH8w+
AEfXwI8pSL/Cl3mruGIhL2F1/PZmnzJWY7CoLFFfTDo0aAfEoQ6D/VRfDnTTXbR8aPdbsrFEE6Yy
sJ2AOOcq61M2ft369TCNDutcORrkNSs3b+UTvuL650z3gyUMyP+zyeNcFl8P+q70C8YvmR0JUFqz
WuWVDVlA/TU6xsTTQLb8v1wULyaTAt7CJ2GrcsUz4Tv6XmsoDHtYHl9mTZdynMwt3Wwap+nyeAlL
B/IR5ugjs4aFHedhTtqeiCnhh2nkM0HwQTA97x/4meCrGzwg7yrslpr49recU2wEU8z2ZrLbUVPP
2rTPY3x+igfaTD2JD9mEotEeV1P3/dg/OtM+ko5Zp5IQEOOyjYGk/cXMb2OUudULUNMdm1ODRBmW
VfYnX0UQ0+YeQdY1ZwG4RuQg+EE/e4nAmavJdBSliZQhdA0xa+nobW6VjkU6VL4CHibrFqCwB1n0
BczW8rfuj/yKgJ9dQXQ5za4N6PhWHjEvR14zgqj6Eerc3BTrf3togjustS9pZis5I+/htnAwntQN
dAOAIoh+yMoAC5LZzp55cRgQ/9GsTy88WrHaLkIWeZytOf02xolNpy9a0Z+66oenJG6CxHVoW1bf
8ZhD6hu8D3iu8z7QBWAzAjVBiD1wZx6/vwAGdIAh2eWyS/FName4d4bWQuLM64HcJr3N+XkFRWrK
eFVCU153F8h9OghnTPyId/l+dAhnSdz37PhS3AcG7KcnbhKLdrjMZQD3zrSxCLlqRFuUx3/T3Aoq
qGOixs+uGl54HkNYC6YbgNR1lNOyuvN+0ZdS4JGBJwMfzFcDgsT5aGKx9aSsi8xPBbhrEiEQUG6m
5kHCpZ3Y+G2PTt3v3ojdFPHrKvTkKKaeROipdRx+JomCkPd9qcueHoG58MizdKzzfwkksiQwGBSs
vOscTp4erXSkwekcZM1Qbr860x/Tve2UfP59Y6H68flII3LzKD7KhoDAj5F2D77YX+0MHZp1mten
uFDmSOy8aw062VMcxtb3PWyATxehHIitR2UwZZ6ETviXWsEAIcmUZcXe9V2jrc/ZsCsMr/a6nJMw
E57KydidT/okBm5qmLqZ5wpMb65cXsDggXyC/tZI+3ev95CVgKaajBwSox+etPsiZXFzbIk/wNBj
h8XU9R32MN1ntWgXjIJEJLx3AhBW0eiie7UiqYY0kJXFDJGVoveWMMQvfxfugOKLNZmp2XWGalAs
/cVoAkHmm22iF2d8m+1jWjVovDesYX36OdC4/ONsemOuIf0+rksE4PtjBDJ76slij8Sb+S9StaaD
SzJTB53objT3BOlvWNx+qO6p8XoFrtBLCoz3wSwDwSsJwKIKO1HE3ZAgrwls9aCxP+6w/r6imXv4
gGet7D/qXBkCE02Vo6koKg3Lp4sZTeEiShI58z3asBd/WNUjMV2oO7P6p7R76ftHJ6wa5dVPcw+P
Qf1Uky9/AuT6Skq1Dj76vKuF0GWNVdcSGNg9N/IEQyaymS2yxIzihrcdnD1ZbGTIk6ZLVfB+Zbcg
8xWJ1eGWRTL9vyIVZQiC7V8vLEAVlM6BQMAuSqpbWkOhsZhi8qNYxpYXA/enA5gHiHQCIugcQI/6
b8/yW3ncfee2Gb535quDspeoBjZpEKJGkmdgRA4iH7t3P/wPxmLpS3oMIy53CMpos/O4hsz3lABB
haShFfBpTA4Ykb/FCCBZzIYrwRsB+vQ5/RzFPQCb4ypaaccQLS+v9hr94hNIf9G4YPYgHv8JyR+b
/ceBu6A5JRNqKjOi9rpafc4L/GyQfS04JuE8fO2Ogf7sy7+FLD2kZg8C31RVOx8WlAkgI/y2xa9a
W0cVgnoc9suGjsKJwv0YcWz/8XrmBxMM9fjal+OezYiCln1MVTBjf/1Eiav5W52G3zNL/fFZzYKS
xtIyDt0NOMMhT4o3lXxhq6rDMtUWZviAyxhG0XgJHZ3cCPyqAUIPHXVG6KW/2f2TsLFKhBVUIm56
t/HjiS7nXo1nVbfo3VWYoVvRIO5iMCAg8N1e9mxBBzi0EmFtiRgLpobqm6D1xgvJLCsNJl1W4C2F
e5MN/bOfDz3v+U8DiTSLY6ffScTn+O2xZCIab2erXunUi6UMc0Kp1HESfDXUijelvIXmmjFX03xn
2ED2/TP921Sb7It/5tJw7lc+3qpnj0v0mt4dWmL4QrPN/b3VmRLRu4YZ9NohGYvGY9mcbyd/e3RF
q4N2L/MRsrr1tvuGOztymo4APsrnTKh0SWuIlW/zF5dTTw/R+L18iENOaJJhPB4jt76QR65MlP8F
JBae4RGwgdpDOxaEqivDLDJr02lsQ0C4aQtsb2qdL23Jexl2c2MvykU7+Y12jgfdLeF1kwtjZWOn
+EaEAKRrLncHhFyjrk2xMlC6ikXCLVCWNJq/9YY7siIolIUymYKa4MkpGDDaoa2hu+GMKsuYnv5y
S1cM5n5uI8ekKXxQ9UmJHiWcGn8TvG3/IrUyz501t+TTgm9bbq7ReF7wP9ElP6FmiW1gW8CgJp5r
DYj7d878ieaQeikNITO195cqWeHRU5quuSOSjzciOWEJfIpAsgTIlfKvTljahVyLd/22/zi8VlKR
jb3gsA8YRftF6XtULK7FG5wxV+4YZizwEw3ZSBSriz2B4NJ9U10+Pi7ZJiM1qaSAD7ODFkPfCyt0
dROnMY7BJYW3LjpMnfSm27tt91TY4SYS0StYJIepzLZPzmztwZdkBMPkmpkY9cjjFISHKwFl9q7a
OhXlp9hYt9ZgRsikXLDKyg0PdP7WIj2ETbwYIomA+0NcQkeJvIQXPophCuXBP7Z2nx3sGdvwd6l2
hg4A18ly8RUhBV0b/rgTLCdHfTKoh2EOUY7EWijPCAg4OrCesq12NeFAs1Taf11xsShcwqANX4LL
SYTAaYwi/0mQ7WkVKez6ZDviBmzedVs+kjYd/w9dBnF9sh747KbPGdFLjrReTvRu/oc7UkBIGC4i
vtI2iwhDpBJBV9adTaptZ52LU038f4oOcOsSLaKG0JZ42MZ581UXz1WYQ1tOmzO1zcLmz2eLoeab
BEKKUPlE7+UCq1yC/sWBu3/Wp+PTN8fCmvzhAHA5ECyrWbJmDXwwXJhyHFO1uxQxTKiNeIG5iqOW
BDdLtEgHwnO2qva+3YOeGyzkmvnu3HymrRMndaKYgUWoM+rQfnoqx483SdwEXVc8M4sgdO3rUIA9
UbAUWjdTKWD3w6jXq07y49kq43KE30+2+Vr2ljUDyhv5purthB1Mbs9XeHQ5aKh217XwfEyLQVGP
yzu6sGbqlbDAuE71RYTFhURPw8ziXd2PxeDxIzegTonYdjNIKOP6lUMBTO9+ooqcNjJmorf7jhez
WY+YTruor6vIaqy4FyHQMnUOQrvOKgiOR02UQM4sK9vRKCBZN6ulBOEWUz7Dtzb/cHIjkn669AsW
dKnr4gQ+fS3ju+fDTX0datflbBRxG5K3+/YLoxg1BuMrBax1D5RzaMgd3CqOxyBzpBRciHlCkQOs
yVVFg/A5jUj5vpS2SYtfTag9OUyOxJYadWYSzQt9czvP9k515MqVP1tuPY/EIAT0GTDqO47YHane
MTUJKs+/lGXKrcHyVtiCl/7qLvqZF96ssXnKl114EPQhqlN0ewuBBy6OL2ASyGf2qBTeJUxWgMKP
QG+0hHYSdjc81trti7x54eNwBvqRfWTioc+eLc0Fgi6KeZPea2zrk8zI5ZBUHv86aplsjjyRCKBB
OGOR6+Y5JoE/Lj8zl3TTdwxQPPSa28rTH0L+993abFJvT43rqnYJC3ITOuS1XhPilibOzXcA2PZy
kPSewPWSLlWihQQb+HfnDa+tFibb6jFRsqjeqWDMQqLGnBoUL525SvXta7ZOy9LMXpKtncl53mH0
wDfYQxKrx+S2CcCtDvjeQDvEfMxnjF8aH6kF+0kUCmKhIS1FzO/B7we96krrfQB1IiJoV97FKz0s
M21ncpqN2+CbFBUnfE1K9sKDASWM8Re4jRG6RheDXx5DrjWwF8NgqEBBCmKrncfuAK1/lstvjWii
NSPaUnTCJ/13Jn9TTMQhhQS/nC1jGWl2iyrepfeLKs21hfU4I/KYMJnQc8Apc2la59UoqXQcIrJx
Bl+ZLjBTzE+ovyLcYFQVvyp+cIhwYa9kSxN9xdTKDoRPfNU3QT/mNl+ZlCRBKzhSywbvmEyVVbsJ
dFSsUnvVgIA5RB9HW71Plm3DNbBWTZ5bdsh08nwqbtllrb/EMSJr3QYz5fFLUVz8typUGGrb8RCF
DlL4Pp54xn7n2aqwagOpNNvO4miqB8TzRbIpov33+Uyz9R+CPHOuA7kVQYtRwnn8Q2qFWA2Z4ko3
LgRZb/ZF/hNe5Q4OE61E3iYB0xELr9ytBrtFuEMwuDlyVxQg3b+EvJigCkXCObglTeumUso2j7Dv
WJIvwg/Fwru9esve2WN13Je/e75E/Rlc2Goervf5o47nAnch7ac8yQtCeS03xqj84gJlWf3wT8UH
a/rVFY+D3D+BzueohSkhFiRZYLlayzske+94TRBV5+tuN9xMba4zVPFkomWLqY4TytpH6C/RDrY/
gcM9MW4dwpiTyWGo3xb6minQ/z2W3vRs4OiclMLrGopO2hV8/MIO0v689srfqPkCSfwlD4D7VN3E
3PdNABQPtv8HL9izOUDHdbKfJ7NelEr/0nQv6g3oReQMTcbFvMfPfVg1YQ7ujMfiCsPkPJJUT527
61x3o/sPW3ylLxDWrv78glKocaeKA0j+hM2lTWhz+uRQu9LxVPGzqwRiKBxbpEgmob49TeKPwMIe
V/pUurAK9I4uJnXy55WFav2Cai3l0yxyED0D6vqtEHWFJnfStIBXSID1mgE7EdUz3wY5IlKEsTRz
O3HaB6Gm4VKlEETUbDQq12ppUfUrQC4/ZEhJVP92LmjeDOCHwE5dNvK4GA1UCW/+NkAWmvSg3ViR
PU08Ukm5ZqRTDGIdb9VQ3evuaeA0xXVO64KELB8yPplKrkZRbN/UF8NMcxLn2fSmtTdVDB30Y3Ct
nY2NzuDQZ1QOEuslsrieEwtnSXHDSHM8NCoCfBvhs2POP8489J4uTxc1t4vzdUPrdMN5SLAxQ0nk
Ao7iEncnuv2KssuElCbVMzupIJr74K3YIBYflqpv7cr6kZdC0+Fs2KUx4in17p4gxDNCpqIlUjOo
IwGSzg518M2UhxSNWLo9zPDcRhsnnXgHExNmhS7FO5WTRz48HDcw8mKow3/KV6EZNNp7hkVicIgc
309KNQZ3mq1NWJW73+D4uRdPKnCKKdnlmZeR59u2qSg/ecB28aGOvlyYi3MvP5hCSVZ1+8Bj+4Gh
LHjzURAqnzo0Il6Jt+bxM4LD2JlcC8NdVBJ7Jj7cKBty5A1peTCRR/v9ufolyI7/85g7J9u6FnwK
hnJCDjEzpRyLxxlUc37OupdfBh4UvpsG+V1pUWBeOl6OqC5qKAFOHyKEi2Pj9dzTLU5ouFgAdZe8
8AvtvCSnTqKAW6lwLzLTvVtQleBcfQahLdeg8Mw0LYn30NUVvujJQWi18WgJJBMtfIuWYYsgEaiG
l80ZtrQnFXgmMfFe9rFuchTIajkglCMQP9vbpQZ2nALaas4qMXES8eSpt6D1LrlEUYlsMhyOchnl
l0ufYabM5XSUKh/H9zFnveGkYEak9SqexiKS6H1LjVf4OOpMjDARbtcL53bPTqzEiaGuD+NsGrNR
A84qoAuA5t+utyNb+nor9LiT+1tUqOImFDz6Bp+okUfhVIpp85XQhE9ipEW3EvCQ5jp55CFesUqq
P0/zggOSX7QSye/rYDSXv20ksIQALZDnouO5+x2/k0WIkGTl6EIj5UD6vEOpC3ARnprkhS53TBOK
/2FC7neSZ/clJzu7dDAkhJOKVCOuMugRDSNIG9U899nsrCOrRA5DQZr64tVCru4suDJMiCOPQ6FC
4UwGq/bw9vHWU/K+zLeve7ipLXUd9ut5KrrE/DBNx+WvculpkM7rgmwhnPqGpUA0z6yZnB/NHmt4
dNyFryHjr55/nb4W3m+FQXJoZVOtCyx46asrOY9P1KzlyFATqSmnrB3jPohfDh5oN0V88XIILG2c
SzuXVM5bzEdf7rv+c/QIEyQhN5ZIcFNqibhuUDkLGURjjjft9psxIDOKUVlMq0ns3xRxjZ8tpzIM
l54Nux0oTX/y0AMgZ34Od/N6J9D0vD+M+O5lNyjpaGDx0C9mYHAbBbxB2UBLzZqktTmN3Smutfvq
7jhV3eF8/zWX6nM2il94bAZHxfDDuB41QnbZZTl0XZJwnfHf4KdxsTk3WA/UY1HkuQMgC9fZtZN9
kD5gux6XUaakY9RMin+/26FZfzX5IxtLZBGlRxLMuwik+JQSaLK5OSG4fmjLYerUSJIFWezPXWOV
VvTDAWEgsip4/6JywkB5TCVBpidO21STFRgE0tZnrC6Cac626cG57vRq0angCoH+neoo8CqbqoIN
/8Tl9pIMYpBhkG2oayQxh6v+o2cIebCQdIWdBhDKV5mFlZLQFteQemmw15Q9wG4w/hCbQDG6sVDV
fnPKdmwmwEBB8XhyQN6qsyUKWPsOJb9awi53oY9qdcZ9Nhl2I2AYHSrtfwRpBYbEMYQOLPYUmgwg
43HaktmrFWFyPRYMn47D+Bpv2wGcLZk/fBNWVWD5ygV7bcQOWG2RVHxFOVgCCCuuN52YBIny1CzI
CB+tTMzdj6Cf1mytTD+aJwp5TDVfWfvB8onLJ1FYNkLjbar5AwcXTeIYBysiDlYQYWVQj64VRMcV
m9lh28nMEaIXSa3wCFqOeeNgiN8/Xu6+O0Ln/PRNtBHIOC8NaVpPS9slrP/XHkdWEW7Pii7xMRqM
/CNqYah+Cc+f3P4bG8MLNoUegBg1FD3KqWSt264kmaTFqeNeoqQsni5JZ38o9v1LPSaFRCcl9pdt
jAbcPfRHggmZlduebCE5Zeeq5ZlMPlQxXcLtvOrDwnSrSKj6HE1t48ji2tyJ7K9AoExAqRgg4ELN
94JFnuI5PQAtDXkP0681N0MxanRlB61w3XTAtmU2N/kzcLYNNUIUqezcOXci2CSrXZcdCNmvp/YJ
jc/NsSEFJUGPvR/80NnU9NZmzLm06vTvbyyBXCxdMNX1gNxdeV/ISXhmY2W5UeQtth4FAVXKfN6N
mPbJXKF4Qw+7b5vhYFQLGLxJQpP6WNOZvR45J/7WH+LsOxyXQaXTMbgQpG2EvA1ozMIyG9/sEQ8Q
rjGVQQUbkuBGlYdlfANx/wT35wa5ek899f0KrVo/xcx/3hN3q1Wpmvz4bSRQ3Q2o1uFLeM6/sV02
l1KZmx6sY+20IgDV+mEIiT2XeXkH+Ecs5SEQrHxOkW5QhamDTYOW2rNv75+IN+rLfbCVThDODDJV
NFDwaJUe65wQR1G6P8lmV9hRDepyPOvLJlfUEpO8BHj03liZgVOilKZII69aENMXKqxPp/uD8wrl
YkpDk7d+sunC3eK+Md5+h6vLClJG/ulRF2q5UaZ4fz0xpHzJgtbxsN54+xFI8jb0BoJrIFwfx15s
vrckIo4Tkp4ivsd5kyQDzppqJQ3yoCtrUNVHHI//EUK4JfDnghHnJx6daXbqd2MexPvsDbV393st
f2gs4RcsflB4XnQjyT5evzx/lAKG/7AqolOgXMHPHmAUtVXY1/fl7YMM8BX7uJVFJ3wb2MnslIS/
PFMX0Qbi5EVxsAJaviN1Sg4pticdsu+Do5LwX1E0C0Wo3b8dSd7o0aApHj/R3PfB2o4d532q0954
q5FfVH/nHUuh4ebjY/o1fpIxeI9BGGPBL+XsGubaQO7LKQU85mZvOT8/pnaImgKMcWBx5ufQVBfa
fhF1DESEDPRss3NkxQJ67FaL8d3ETWb7BzbwfHTFsuuTJfM6sbXAGRYeK6VnXIgvmwMteCsjaYBy
xDep4IauMfNYTi4ziMd8pKJWDS7cEQaUYBjT2oKzjmzKcrPQnLnrOc5YNpaU8TMfBu3DkSzeNcLS
nLRTfZ1/6OpUDrKNh+Rm6wDQnMmpGxSQj000rQTDj5suirY4Q5faYpY4YpxwpHgTzhBqJoUYd4ZF
OpX9LySKq6iLUa3Z78DQvrXn0+kXf3Opkx/ZNoSOd7Cmli/qItLKQ4UNRNkO4hno962ZAfo3uCQP
gOPPzFxnKoDOeGrXbLqZQ/nzBBPu1BNJWwpMJIJcxxy33fr5LLKO77TBkqH09Hbv+/PyVWO0U5Ky
vmvwf1+DWV+9ApdbSp9eB4QpbLL4hFrpa07+bEHWJx2/cTDtr5kUehE3sEHZX3Eo10MXI3SMdtWQ
jMSEPiNv3AqxdNeUNqnbLC1VUAq9CpvwQymjOu1J5QMz7S/oGiOt1b2MQyLnmouWCmlH+e2m6jgj
a0UreDe5OFy7jXtUyI80ZRHT4MjBffHrEVqa/zfOpkHds4atJvhsE0PuantKapi6tUrKtNsbyVJG
FXYzwzdgkolJoJhVeCI002tCACcbrs9PjsMx1vc2sxv+aYjI4D+WYT1K8JpTj08eOZXuMieGD38+
BCUQZLfXDTtJlVMqOzXK6rBbDo3pGnClsulafcuXWm4IiFdsGZXcHcAWJpg9GOnGkSHoFEVGIUcn
VCq8sfqVkR7MYM0d0MoSF1VkbZMGyusDnl7T7TVSFHbGwxPKnPGtPJgoLnJqrtKYtAFrI5xKtN7P
4P6V+GEQ3bGD7hfltYVhXptO7I4nE8veoa2dKrlxSoO3Q1qKdWYzW/7eYAjDddkvHGNxr3IYSd1N
VTZ3NnvSawVEv31Ryq78Mk0IdjPIqM4UGusKDBiBmWd9lGcYZg9HQOnOKLPSfTKHgu6O+wuk77jw
vvIvV5xjq0sV+V2iT6g6f7Xf0E/S3QdLg8+cn2hwEqKsD9OzYPWFKjwkEaa+YSRU/Fax6P5jUdVI
Le/sulDpQsbqAXM3LHb/4k71smdU3KIEgw/rRWaMpcAbn50yZhbtUQz6Q4VT01X6CYZZpfxAJIFu
xTZ1rmH96XTPtyN08gSFje+Gn9YWh2lLLfdDHoeR+J4ShL0iVZe19/kipd0/NVb0/nZyvapMZC9p
Zw/YhOL2AXMiMOfc/hD0knyeq0uOh5JG0C+COJmRK6SxOJGKJKOqbHdLcEl7KfhfekIpNzFYL18u
F7Q3jkheil4S9TYg6C1TnN2Nq4NwjVHCr52l+mLa6FZ8dL/7h4y+uTFmCes5tnUlXbnQij/JOoVI
YmjUmDZYj5VMG/N1zS3i7a5H4O4MfyAuHT0MMFII5t2tSW3A9Q13ZNWK3ZBFWJlJppCitB/8fsod
PPIp9IEPmsiFX8u9qAjaJcO0jRIYDkmQ0SdEH+5YM8m61LprKN7L3c8Yku/jXyBVQUJdpI/ZOfh4
183gaYOOzi9WLjlrfejv+6/KWHT7Rk458zVUmHdT1SBZq6646ZmP/N+AVx4Z5v+Tn2//XKAV+Bun
TJJmuUkTF2DO/GP2tmVlwzyU0icDwiIjNWARVvxl69tLQpBoJFEhTQ3cwT5lZ6LZQmpAVkACbeR4
PSZubxCI2X7h42ZrqGSBDkzaICiyraBMsWgApCvlyGVTxJdgSbMztsz3wG1JKZWgNZnXqDt7aBYA
CHttRx95w12quSuA1NumL+HA4AxapndBX0qKjykLEbRLX3AdGoYIWTjmtrXOZ1RlVdDCcQI3e3nI
YjD8u101xzAJYG4g3bNdxV8f567hi9mY900vy1BJwaVl8g4R28wtjCojW+MOJdanoYIaTrWcvb/g
Wd2NIQ125L91FneMbXgfeUVpES0jc3kQwBZTL7p5386x3s229NtIFyuAEGiL3WBw7GmQ6s4HdybM
H0KJVS2z3Q0QIqrfqwAqUqFTS3myo25aPy7W/fUQbqsHGpBHwt956/8IoLq9ugQEkdcBLPVZqWwQ
CnlCLLxt5eI2Kz7YA6N9jO1W0eYs4qdoA8qKGTcydWAZ9k209Xgw7PM1XB3U7vcTfMCWoHiie+hb
uqrg1rizoYhH3JKDayLtKwk/O88PtoYXTLnLXkmLT1ZfpVn5FOgFAVvaH/awo2kb0fwSdJtOETc4
mwxJGA4lmKZxMMNsCVNreVek1wJzmdGno1xh1pK3+cvifytHKrQkHM/Z6XJGkNi9H1vNoHDER97v
nxMPdKWc+wcLD9Esuf63vr4baVbFl+7BRGedtPxbiWbJf33tBOBlSl4bW0stWFfejr+aMSG4ituR
cPWN54vApg/S/KDREYksDI3WldbLqFqg78MyCfwTBxUACYy7o3W37QXFMlq8qQlI3I8i2OTbR6Rp
PQEs0cDnLbbF0Q94xJys1wUo2Ztbawek0S6GTULW1fT48z4uYUvDrQvz5A3X+WUg8UwLf5Qd+Sbt
qrycLZpWCZx0uqJLD+1oCoRMJW36RBRnty0b8npKbyqL3G22m625HkL7ag8Lq5yrUjNd197Fri77
Nq3it42a9Vu9l9/mICeqDp91goTIZ4mYD5HFSrL5OeTQmVvSLANdNu1P6HuNRllVeixBkW3VEcEH
KGOZW2x3cHjiXa9o8XaMjkNHxOU8Ahmvh0blZd8TeLfpXkzutf0ZGZt34tzducUnc7sy9toNeuW0
Zdu6zxM0mFbQgAPouohUnE4SU5a4HDGBxDFGg9rANgEDJ62zRJw3Bv9G/W95h3WgUoGW3x7UcgDs
M3wHrF3rFIV+Q+MF88q+HUhjdPIZIChnxl/OFYHhEIPXae1E9RgQINucOLYqzeWnpm0KNcV38y4A
3djIWefQg5gaHUAr6yJW572RM1+jxq4Ytwh0zVcXRHu8Nzq6RfHxW6EeFma7m0J5jfI3+bh1xcab
tlHQdHrNh09Sihk1IU4rq+fQhtOznjpZrnmmvfAcTuXYhSIkAU6q5e5pi9ThgkJ1rV62msz8uFQK
vFgg59/MUPRYqhhstTgn5soMkyVyKh0bvkZZUmWNwVzBy1bfU9eZ5XA2Y/oXWSSsw4X8E/rNgJTx
58B3EDmBH85P1rd7dTM/GZgI/gm4nR8wOKFVfVE+xSjmWcrO3wOl/04+kdhFWbTeSIqe8kRcBUc+
L8R5lMcDbx9pzXz8DJwtxk0aBRZdZKRuq6Uxaacoh3Qc1WrdXCaJSSMUA9N9ZvGbLuUhj0Eo1sMD
WTRBd6+rtVhRWzO0oJg9vfN3eR+lXIXbovj0Xa70XJem+1rEY0vtJo8rGciqqe1vrvoGey9RU6Nk
722/917HDX6LO7+pGWmYddc+rFhO926dvhwjjJDOgRJdM1XlzIVHpdvXkOpwzjPvdyOlUl8aSK19
Y6+XaNTD9gpHSy86XZU0JVav8mzCtRRIubr7Q5PJG29inaJTnGLkPPIGByxiMsgfvJr6dp6y+RJY
yOvqNh86F+fLhkVFRe7NQhynUmFyRAHUJDt4jAybx9TTYF6wf3rApgaJskxcGetT5VsfLTX2+g61
BjvAUPk0eN8ySnGWlztbNROnKECWpVW2PZlMbZzanCVU9qDVlLnxvf3o8cwqBgpigmdaPULM63QX
23/VU3OGf2naojtJSqh4saB/wmMKIYN1MT5RFEFGg1alL7SrsU629QMx3Sw5gqWmG4EMs4JY/vz/
0uTcd7V+jFvhEmKUkRRoHs0QCv1mmPU/PugFQPONpjaVSWUrdDWxLgsFmbaXcyMZsgx3a6sJzC3L
oN186hdwKu/IVMmIGb168jKyAjQBGuwzwSjx5xSE1GforrROMw/6NT4xcyJMirssVu4DSHEAQP2j
pt43JpO7MPdFRYjp2duLyzWz6NGl1PKZEhzB44A6Vcy4GxM9lB2+142+8ZbUx7LLPo+e3YzJlmJp
Oa3+qkKaRWMYc/XwifRPFjePpLLjc3s82is4bJJJj08hvD+LaQSJD+wAUvxbw8j/8oT/ntJuqGuA
Ermt/hVXVODvWIcC/sSSlhJvhG25p51kB4lE/t3wuAINmYBvGsjLR1h9gDq4ZXVZzbEJcIW+eJEK
0iA38VLlyPf95AP1xE4dVNV1XCkRUieugZes+Lfx5U4F29eOsgmO4gfMVqGrYV1njb/BlNIbvmFz
UBjV6vpIyPh/u0trv7eT8bXQnSQnJkmgeVKxSyE/uYKH+v8T7IMFlgX9bwyQ1LP0FdikZSeVyDpI
PRj2u6daqfLoTAmfTcW+Wg+ZjT3t+R7/wFhchN/hwkWsZY4Yq9zrGbwGaGt8eVZ5dIA2uU/wWDEv
RvqO0dMDwFiAxmTYlMYkirl4LAR3xqFH7q5webn/v97I0v0RTzaGvp4upUeukXDrtakD+EmCS9/q
VDG/vo8c3sbm5+QSv3dAjAmbIvLguRmGfaGZRzYsrGqd7k36HY9hjWj/glA94U3Vj+jB8yE2of43
cFJTJkOtHz6TkAJp+n5pMsORLMxg+LFI5LlKPrcLVdHiSFO3YVRq0MK9nrcAK37PQc0adZkotTPW
MqSPraPukF/0DSa1xhg42fAzVYuzM7bTo8eZJ1rqbNOAU4KbDCgDzHIU3ujqBDtmALaM4C/Ar8Tm
6aRTuS/qLgU1dME91x4jvX9q2J3RJcuNdGV68o+LsZvjSiBx+LLKxk+yebNKlUkYh/JiwFKNQGWf
PRKMs7R00Y8u8DShP6TeP8uLTJDs+jO4IT9o+svx1XyaBgELabJAofw16gqMJugJ53iqyP1C4lRs
D8vtPGd7fgKz7b3U11Bubf+veW6GGAKQ4o2RUHYC3C4E43FQtmOYIAFCdLLVx6dPmPui58x3ccB1
cUj8OWVfAeOlHavMOHEHWpkDXcCMEb9ne9K/wS8rM5Tj1ya7LqBc+vR3qqDmpaFWGhVATnHzYp68
SU80zq/5Q5osb/UJLsKaSmZtlWMyt59oGLGMqaL3xaoSg0N76fGx1v4/90bF0JGJpW4MJgEIT1U1
Elf+C1F/3w91eSjolzvVDgktpECsACmRu/Ct26vC2p7zj/4tRbm3xWz/S5ucTIXgdL7u7zyzFrMO
LItqwN7X+fch/SouV51wTjsmVJaaH9k6DiMim/hmLUpUn48NUiBBrcOyzZKfJzCDmHO9JJIBmIdl
S9XIJZZfoC0kKB/iQzFb2rXDWKDduW8h2arQery30IodlT59v9xFLNbrFil95THbb3hR9hTGEb1l
y91Y+P1hsVON5T7o1VVfLqtU1DqiSK4VspZI3ZosAXEWGGglmmSFdXlwEsS0E4U4lNIH9mhVy072
uVNCr76JbWBDi1hc1r13i0YXozgHU6+HZY2XWC4AW7iMvOddoCfTlGzvSJ6yM9STeK/PcrTxOHFD
Loq6XBMiBsGeddDvVTugGI1EVNytZRWF/xBZt1e2IcFmFkloNAOfHVOh0+ltxB2u27dGksrZO17P
2yl0tuvvp2vYjbGmxjI48x+1E0oghA4z8ikMEkR4oZSixSAInQ0tZ7lkGREfyZOGnrBU++ZYwYE5
ybhHr32OveSlh/x8Rh2XKgzVt6T2z4jHwPpfoyi1lEQM9X/ovpUZ0NgfeUJwtBUPyDCi35hCxlQP
PUXL/fDNjPMNSuJgmtNqhXcSiaVL+fed0UBp0EOPjaeH1hKS8B+lu8VKdiSxaq6pVV3VojCUplbj
DX3IByWEEmVMl5j6KCFxHzqyiZW58Y7L+9FFQpvK7x7JeUWU5HOJQDKqOlLqSMr31s5kC5PVMt0t
6KO+RkIRDZ61i6+NznwLZ+bRIUts7A5h7HS7YHKymUy+9TUDlq+f5gNAEhgofnYCv7oKaSbGu8ap
RdHiL65sQruPnwtbFR4RTplnfqz8GAnX8VnhDolF1dpn9r56kBQ9KrhiBgNvhTnKC02wRPaHGrEE
XR2hr1AbypmgbCwDhYhKSh6MEPp85xWLDqoXAyqtyHCCYvYkzIRESoeksj0BOARz1Cqbtmqz5vHS
9CqSzs55ROTzE9BRyWNi+NlNGvxq2IN76zROVVpblP7L3qO7PskXbsTq2BBAQyk6Zg4eH13JAs62
K7WwsldV5MFgzoZaMkzjHO8SMDwSEfjP1EjOzuCgpFV/Wi31NfMfLIgZ1LKX32YC1JmmFQZdzVzp
1bEwuS0Aed7QmcT2hxeLAQYKw5IapsssdcJPrK7OjxI5y+5kQmQH5UxUt1+i1Boe+Lla6pHdgPVL
niw3nZh2AR5z1iiuHnm67cTkmtxD/miy19NhT3gmPV4JyhQQl9PeYGg47F0zBdHMgSOQ33CGQ2nB
CvdPubvnYVbgRVAVM+z0BXQ0mqqJsWeAhljzYvRkHKiluBGGFPs/h55JFUm5FEGNE/hESPZz5SjM
cfHvFRRQdEW3dRnD1vMfc4jUFI/srcXsETRX406oO8t91L0RH0Cj79l07hBWsdr6GuAGDpD8aSa1
IPxPr3H0U2S1CM6I8AGGVlzhFL/+GU0kkFrRp/oiAJHZd4ecegAL7/gtQsSrqfgK087gdrwBuBKW
wiMcl6vZ/hwdpwYTZ0+TMwyCdP28+LhoDNhl4GhjD4mwXXI0uRiBr2cBFxPHxB6WhTujgGVN6uQg
V+6/CpU2E1I3TyE7IBKsuM20D7OCbfuLpD69klMHzcOMiGs/X0ydDPCGkiXYaAVbotey5klZPJVP
C2CQZOh0pFBeCzhPhehDrUYtuOw5YT/fSYikDO0XfhlgBwyVTbHs/EGM8zY7qA3tsZCLN0JFmyvH
Rv7hHSs7K06Ct/DJRgMFs6VxMKR54T3iQazoOHD2WKs01jN1hmYLc36PvXXm8pa/OyHIVGLiLjQc
QbG0NPmdnIvQB2u2cXRe9M/oHvE0JGlXxOxsI4kecloQzY6rJf+xkDveE4TEvLA3IeCQt8YMyt6t
LbFbXrs4DhYt0tgW5T6QZU97MMo0y8WuCjUqlauxszMkdfVJcUSIVIFaFKfOSVixzkVPLM4Dmc4t
2kP08CcEI/kCDNZYLjRoJR3Larh8nocnybdIc+si265Y0gOJP1Z9VNKlXocKHfGO+UT15U4Q+GKE
HvHEO9vI+V5gB8iEQkc+BYhuOQGUkEmyp/cs6NLfv3JndUns0PQDQs9Pw4uy/OOCB4f+PvWPTSEj
xZHJdH25Wz7SQAxdXSaI+NZaz8mY/BFkLCQUoWthQHNILk4fJQegHGrFVSBFIV83ysfELIZJOejk
NY6XJaD7CgfGxrpRgVVUXid7btn/YehhhBPoUB39IQcd5Zds1MF2kOishvJb8JGD4FaIoUckaheC
xmAwA8CLIDsJTDuy/2KU3cTk200bgf9f/xwIW9F+NpZ3SOM/+L7If4C6N9FZ5k6Mmt6xtwSRExvu
1O1XzkcnkR1uD9D4XnPDHm2XUJvaJFLAKJUoPliG4zne47I53b/JQ983R+CIw/WwuEuNuQeivWhh
DBMzeX7nIpN+BXN0w2dAaqzc5qjBty/lhiAMLohWGgkmewRy8aQ48ttjd2TJUUSIS8jbNoMZLEeG
4RNfsEMC2cVPwWrN3XdH2PrbYYs3JcIRGQdog/ucwPrFiTRYQkOZbz3b1JvmrfhGP7mztWAQn5ar
CWnm4A/kRBGqZSzJByUvPmQGpLcyinSgSo+l00+johHOQAnFrg+XsRAPIMOMgQkjHEl6s66fPa68
I/fl1rlaE32l2/wBoymD/4gb6q4NVo9GXkHTLndpAgYIBTJhvIt1jdZwV1ctm2DBFEYbDOdnfcD7
+o39x2oBXNhGj9tpbrWGruVWTwLPZnVviPpalqA0Ex+mV9isPCZjq2JV2HRYLjU17tQ5F1861cW0
4f5EcVFRyDfNCGaCTw5v9lGOKw49F1zHgdcmRABLOx1sceNBbsnGO+GT39mnOSi+Ocy71M4X7Mla
w2GdjSdCqfo3zsvdtj2gTUJE+cbAnglY0sy/jcWZ6jb1t8OSNG9zPfIjE7bTg5AEmvWsyz4UcMFf
TEVCfkD+v2lRG9ZipUpl9pp/E4CVRpb0FXtJq9mFUSVhMl6OpHN1sPKUe29PwSTt5oNkwB0Zh6zp
Fjv3mlCW8ZM4MWLEa+7dYRedWoN9TStQ97zP7+iICG2NqTi3zEdwyvtNXTLABGxY2PIzBAyrJZ0U
HKaIc0J1umTMVuuxLaXMp7hFxr2JViqml6SNHxfq6gcpsNc5u+iA1Bqx/7FAu1P3PBlwdY2hBEFL
OCApJ0v6INq47QdwKATDVdfCD1H4CRwOnIDOdXQamS23LBL4MyAy2NsDPLyHZmzVmSChHKRR190R
ACYQV0hIu0XFJPDKs3/X0d44Y7xS0wHopnnOa16GS0V3c6UnZC3gKC7N1dErcfcybQmoh6nno8DE
FF6YfeVUHm6MxfS5KdzIhxnRunSAAMB+LNpQfDCiFsWLNerr1VRKEBcQTWKI7xLIAFFaOxSY7+tw
iL2jx0yfbjD5bE7ABD+cEen/pGQFxk1WsyJ+DZovs/Gm29R1lzuZGpXivPrG/o5U3UFDpIpDxS1A
rF6ktoagk/YQXNDZ6CA+aGQVaDVSearmRLxYZj3uI0QJkri5eF0Stdr4p1vGsb9ycj+BT/NuP9uq
N8QtdOrS3AiNgFHpkPhhegATC7xK8DSIdGgN32SUS0kRZW3uoDLZs5D13PxmRLWQOvhoR1SwAQ9l
fhsbk7WPflazIvWMA7sP8yJJw/3ttBwYiRSwWCFSC7OP8qYIoGyeFxkhLJ6V142OE8R3TS2tbXJF
z9WrmDVHhYMWv8hxxs1nsHb4I8Uy89sUaKj4a6Pk7sFj3k2QDC6x8ki1+HAPDJIbr6Y8J0TrF+UZ
lJUGKrzM+XPdzVVOpKaXiPZyxCDosN2ZUhPuz6fOMl0vc+gdWCQkE5uekBDV7vrzC/SsYDRI5vea
3U1UbNxezFnxALyAxTSoDsNxrVWIlQ7c8QQyg4VoP8M2DKMv1Dw3nMyuKbFtDh7rZOqUS2qwXiHq
hpvv4xemlCWae8cyPU3mjPF4CMZU+BqMC6eiFXekzO4TjCWCS5CWV87fx83Lx1TKn76DybqJEdmG
eOBIHDBuQXEgUwtCbBbfh/6kbkPME7SyZm4J7yHGGgyMQuuM1DEnMTj/Ne9Yj8u05QKZWLZQJlpf
gTSwipIgV3zomzlT84mbXQHQRH2o2dPyUsP9W+UJOTb+4UZKrreto1PqfYJnbXw9bTDzOxh1DYy7
tO4qX66+PuxjcJX18w2dTWQklfD0hrg+cqq4rzoxrBIT/8plM/Vb0IbwCP4SRPDMCrp8wN/C030u
90Aw7gn9ZcLRF3JndAugrCuMk6AAJYFaPdGQMbsdsphc5Tc1i2QYD4U4UhgJGk60ePAoe0rXlBRS
aAF7Rg1sN2ZllzySrxwEO4N02jTus93qkNyIQ3sq5FnJubBi/iWBX3MpI2RiikRiU3x5Dxkiy/O2
rYPOiBinMPMy6FkYnBADDOxNTveo/5xdeZYFtwoFVTgfsjzTiAzc6kk4tyQojmHHagDNtcI7onKO
NU3MgWLM7rD5Gvebmv/FH5V2NwPzfCo3eEhJkOEhH0KwT1OaTDjPhbRC4THQb3oScz/ICYmjNmPl
ZABZpZTW3wNy8z24j1SbSp/JBk2t11vNieqxVnbvZPKL9lBstwsAH/TjWyBGiaJLmjd+u8+wsg4h
nTfwd5o1oSQ1qw1Sqk5ClcyF2ISv6z7wmxseZeO+27LQpzbJdP+3z+2PL9dkZO9Vg/hKRnz4pWY5
iL4RkjDrV6QKN0fT7M34bmkCnjOY/HEBr53JgBN0qxnLD7nwdrWhvROt3wInRVWwkNJzdM7W1P+C
ZrDYoufSpAHCo9DKoukwBw/5SNYzOl+v1OPGCTn4tVa4ANFIttvwYne+foXPGeCv/RE9iYPXbhyp
ELOGNuiiPOAGJUDS+g0JcuctCSb0pRA68OohocnZ+OsIVZIcUSCaOakA3XnOiaonuCd1pU1zsJmw
3sYi8AeKzbAFxAFEEZLoeZXxDDpETkS0SDWLpNglOodOjKEOJ0o/h0Kr8dXHU651+WYf/Ab7d79x
1pvCfbh9wyUkf1WbU98kw2DcHNpqsyHnzkSzcxoBI8tfn+nS72XqoF/YmcPLlORaJPrzRE9TP84P
10NnXK44okPMrzaU1BVpNIGKMHvcBnbdkjlbgoOZSvjvH2btxMC5B3wRf4CJUQD9NWEBmGxChceY
3GS/T3tX+MF/GVIUkb8wDQbG/u2VZlgdNepWvdiPVELVoAgHUYmT8E3oJS2MtAk1PPnmcTVJUUJF
Zoj8haLNmpGfaqoWWzrGPF20qoAYJTgltWjCUbDjI23aT07fHV0hsFi3hDOGpJ1NxjQrXWnR74S9
eiRh7XQo/avFvFN0mWID+H97n/BGoz2muMruXCdX1sUVnR70jXrgKUyN+vUkUv/lfLPMzA9UWUgR
h4/LNcbe9pIjIrk6v794P5MjuoMcEtJrHLeYJHIwjPYsOk87XFpEvtJfVlTNBne6/alYTQNPVmZl
jMy6CGecBy+tOQbJ5oc6Cau/C4o8r2oK9R1SmZbOlVac/TKl7hi1f1WsM28UZtaDSfwxhV9n9wxF
nV2cy/3i5H9GvrM5jwkP+6d6Y3UDQbluoJhQ/g/rgqhEr7+qzMBBUef7qKYKLN9OLwwiVIQK2rT8
m0Wwx1CXey1QVAn3mFd7a5uCJlaTpzg3OWueLixZYa7qX1aTxciu1cFT0dbaoJmcmQLhmiwzXgm3
A9zIK7l+sOUn+YAwK+youxqdD9IvVbu5Zm45KXhGMtqZ2GpqeXrpF6mVjX2yyvlQfoB/mtCMVvbt
n71Zuo8f6xL469UOIKbvLmEJQnW3Rmb8hfkSAyWeeym/EUbmOXHuKTQqxtHc0EXdZoAC8Soy1o8r
9nJmGioD603lPvUYRsDwsXp+Kyo1rJo5nBlJTXC4C/WWA36/FpOgLeku7gp3yf0tbyc2oBlWs+jV
h5g8sJ04PZUstfq8Gf5FUp6uUMbOj2j7uWfGT6UnslM77U//ST+RQaizz5uuHq9AHTgKWMToZBKc
WnAci+lxMAyGP1T/b9J5y3uXhgDEQZqQbiBmtpz8Qtwd4t/ftxh/4hhtiqe5k4EAzLT3raebKaZN
yH90eS8CR0pisvNK1MA4sdMmdFfq1acUK1WNq32OFF7ypXDrVRkSOQDU03WARQC1a5jLYCx1hSpl
G7Qove0tGcCortLKe9vt8xn/NEbWcaZkYeuqnUyGMxg4aw79AK7+9lOBUsFLlzihAUKXvxw0Yl9D
lIICt7Qi8Q5pCBaXENSWRBdq6h/u73uJVTa8f9tYv+LgW2FOhHc/fi5tCD2cHucPiFOSdZa8UWyI
1lUpre41Kw1tuQOETTKwZzGt2d5oDU7xqVdvRATzH5eDp6IFCSxxSNPaLp6AQ81PboycGI8aeHkF
2n21Hh55Z7GNNIlsXB1vEz5GFS25I8EIeCYb6h56gdAGKGoSAtWxv/Bc/eyBPmXyK1vjkV+HSp+x
AKchHgyv3EWoK4hc9WvVylj0B97rF8QHfNby0+THt1iHfgEGwS11Fr3mfgmU+xHvAj6su8bGZ7N6
y3nW/ZzyHBN2rIGSsIBhdMKg+DWSefRNJMns1KRjoJbnaWXkHKKSgAcTQkW22F8ABIb89Voz7Y7A
gbTs88gj0IH8BIJOKjBsWwxSRAEMtwEeq92ams1T8Kt0RTuWNw5U9ESmJRrXgjZToAxd6Y/ryLSy
y56AbbrFHj79oOuFzdagbpnUR+yWoBi8O5k0Ict4fgvXwrqLS6azTxXcWjDHqKSgbJddOdDsFyd0
JM043Ep0ouXxrHAJ60mjbWF42EIK2a1aR7wYXS/tiN6dN0u3mrtHCwwxHxZSNvydTlVuyd5rpBqI
TjsUK94e/8NAGuKzcPw/ZM4Mh1RmWYrnb59lo4bbcU29NDdm/BZnEwI0tP3e7Z7ubCuiAsKI7L3o
mdF1oRZoezJPQaiFKuNKQGPjWLuXhupu33j2G4VA55f6tlYyZyBqn9N3pAgCo1jacfQVPnAI6eTr
0do2yVQTKaGybnjGQN3vOMUU0YroWLVxOaQsjMIn1MoXMccsxu1s/ze0d0tjd4q78N1ZYz/kCRZp
oBNXgOTP1jCcjq437Bhf+kjD+WpfSAtBj6R2tcWe6SoilnIcfBuuQzmpPe4BNyi2u78Fh0cv/yAg
wVQ5xl6dYgUys7cGhsCQKMl4s96oJm/e4nzL0b/uOh9+/Vld/xKmUH2oRXwJDXTcKQcaZ5cJa4ft
Y5glvlu/h0xb5ezGaI+XivaTJOE5j4WwtNNb1jaxfvVUF1aUdMkH0pb445Z5ianfGtzX7X0T3ceR
qvw7+DINEE+bKc86DTlLBxr8UrnTnETVrw2aWs6Q5Gw6dN6jBIVGmNK5VTiLLACFZ4e1k50lCHU/
kbCjVUrHhBlfUWe3Otv/D42VKAbLawXoo4tB4dKgM0iobjyPUeYJbHS2ZYe2/b/g2VXlHX6sHA5A
871ohxWIzTZBZ93iFqzptRSuU2R1owIQBe37xiAffo4CP92WJ2lvzVKftpIcyP+MwTbO5W0hm3jm
P6HujcQ4U5I/mPtM3vZ4At5uFKSgI605wfmJsGe2pw+ezOb6oqj6fTtqs1080DNqySImddoA1A61
SIvsVddf+o+yEEjL5XdDWOUuoTqekYn/uhk1xahW3oVE56qBk9N46qW0DXWg0ry/SWWVvAhYYOs7
7srZYopSxE8pWAvZRuvZfl8eFhmzADfH4J1n7Lie+0g1qg6CU2cWH4841VXIOxH8TZoVziCfn8K+
kvC1oI8QbnLd/TFKw8oKb4D4I4REeeRQoQ9SeLFNo8b1BbD97arCjYyErbQX6A5TZQxg7TLByM0X
t9lRXHsb0NZAtzmXixZNkix4d2DETSHAYHok4iMIiwJpOen14mhOETdsG+sVZXCjuoQ0VnDNfe3d
Uyfdk8w+9MXXswD56GTJfraTg0KincBufYvcqn/cNRem5XD9FJv7ftHlrRAZJ0IrAAld+tP2M0FR
7rkOSWmPT4hoq8xfIm8SywAEa3yTf/qs7gLY8djTNcC8zZ8KeG4hZy8IefpS4jQco6j0jYWUfMMp
/CyiRdyYAV+4gHDMTZi4Te6KCVbj9opgsFD3f+sgycloavxjcVxOIExO/gyL9CCg1ZLMQhypWdoC
oSNcrL0iMavzc8BI23F92OgTZUS3wg52dYsplC4alKmW/npfSiRuHLmG4RxJe2VyQUPk4JbrOhVq
UDZKOtvCeCKZmTbyP3+SySNsNzQAEjm6Bdp0sfPVEXT8DEnLFM3RDRAT6RZ4o6ddPqAN8bFPhD0j
nIC73QDkE4WDvQSyKlJhjMWTCNOOd/qpDM+DhRpYQYpwEvabFR3mPag7+lmskCbClbFN/JMxt7HN
h1V91aAh+UxE5zNQMj1gqeZ0pr7yNnz1uFDyjCQK4GY0oWJiJ4oqj1hJj5wB/7m21k7RPz/DS9Ea
TaAYOLFQfUu9jLaNND+/Atj5nU6cx4tJecIchNsiJg76oBdHVQHO9eBxKNcnZeTy+1Dy5NnCIDZ/
Gc1Moa8flAmexZEwsoBp26A7lHk2WZICe912BPn5yjt0U1L+uC0xK0Xdspk7HjocYhNA4hHTVwes
ImMn9r0ZqdheHGx9H4HaX1wvbdPjHSGBdqPeoSquH76WplfOl932fdID6crcGzK/5z/hRmTfTa68
md3hZITFr0y0A3tZBJKE1hJ+21kpGesdnuDOiHiyl/lEegv8kivk3+LxzUla0Y2K6gFKmfub8/VA
Hh1sRHTVVMt6MIPO2TnWrue3O2B/iicN3BfSCSaB7sWL1vkzQO6PNEOH6Nbc3wCTsG41FRT65yYG
Jle8ZxfPlotiDW7zoJsj+z/elzMOzYK4gSwXhEsVV13yzQISAyP1+xNTtflNeGi+I1OdOvAKC1tv
UbQNsKlKhDhMLqhOUA7uRvm8hNJy/lO5KpZaSQY3xcEcWToluFMyKFOCfNsNVW+zzMXfik1c34f9
Plix6X4AggsRbCG3eIUtRaStHcZhS8ROfxJo7shcA14xZRU0WPhq0BIU4tkYtrMHx5nCTdAPGhEj
prbewcTPJ/L86JgOQpnM4QZxiwYNnxSsMZm2xsSP41ygtfG6FGWImBzF2Crm4faXkB8UmI1Fd3bp
f9UJ3ohIJFpE2fK4AV7Efcxo4tnK3hBAO4vg1xuTraPnUxn+wsHE5sF0+Kef8OCgPhhmPUBtUC2e
PFt1lOMXX+u+vo3psaF7MJE/R1gAV5H2VXSPuLjCVMGpZzLAfB0qxE6VzjukqU/hHQg/apjWcPe5
IVzTCD+stjUKKan+P5lw1/c2l282SQPweVdbJoUoUSHMDqvAc+D2WCBMowFdnpvMsQGh4i9prJkt
c2LmZoqH7/uceGJFntnfS/0h9/hDa+CYqjy/cBNHvHssbq8gF/4Bm23hx9ny3CAow1NcAtDLQyin
q62t9Si3jTcd/6qF90DHA564u1z+1BnWpcN7BfbPZplRMKlAptehZwRcVxw0HRsgvH61XWO1eraZ
+YhXsWhUYKE/QtdTsIxOjf3qAg984FGCPrSo5+65v+urdUi6H3GBv+YVkCJ/w+hko2bJmnjvr+cn
yzeZeo1p23Q/hsDV6A9JHjnreUWZP5KTtXkgJgEwP1unGXtpvYlyKtXO5aAGtEVnGL8tVdkCRGDc
GQ8yAHh+rie10NlShAMp6QUF4h/xLd4WyNuNedvUqWbfT9sly5W5Fh6zAycPsrcIIo9dYbWZ1QwQ
Qu3St9d5bBJrM5b87uP814HOOYi2C49n2CTBxg/GKkxVh+Ic+TJUG6L5sOYbfJjj1n02R4rTQyVi
o8fz1ruIBOUn6pxDEDOED0ebXLLiCKr5EA49gYVmYbXyqtM3TbSOfeJNjyo072mc/hfLr9Clca2n
HfvJjHeWT3R2vjc7GK9ogZ/incEP9d4h7IqRqQopFPxgSNDu/ohCi3p3MenYgIuMOYzo9rGHACVO
qVTa0a6cPciBoA31CCFXhgQpVqLrxpZY8D2HEieK/kv1V1RiItpSJmLDnteHtyp7+E0dbBULO1dC
YMI9xQUo6lLGhbA1StMM+EhA5jYqZ3g2ksph2ge/M5cGPzWiJauHjoDykdaPq+TZQNQCoyNeMH3u
52MjeEEqOEYoIHKmm1AFfeMvHjTF8BA9aVtQCOpflM4QmE3ORaLoUtlgn+PeIc0CjKcnpDulkuy6
9Toc3sLxgcKMgBkDeGDJK1CfL0FA7+yL9zjp+4RJl/zLPLAz9meKweBs2yZfJvSvigb51kNR5Vx7
WYQVeHtMDaXwzoAwCVLNrxV4VyZ6GFIYV4eKHOQ/4JHh/AuWc7a7sGTjWLjoHSz7/1Ogy07Fu6rp
MZZd+oetD1a7dbedZGcGj/pCylpHBlFjUSbqlwuIhIa86TlPM1WQuQC0N8LXCnPXv4OR8SbCoPQ0
eDFGs6k0XolYrstl1d8qB5c2b4wTZNjSe9O8ZvTOWG753uo6UQgq0EdzcOY2VcgLIMotFQy0u7Ya
VtIs1qSDlFshpxY+lqHxj6j+Kk+Nn1+qsaDV6HrCjxNf2boGr45mMjkonu3PSytFh+MlNCa3D9FM
cena2q/8xcyVigDH/17XPgd29frEP8+Pm0jYinVaWyr7aoJqHYnAzjPo+9wZQKaYm0qPGKAjdfZD
Z/LThlTSyeEjvPPRzvlGT8ICJYO04hmz7wZjx5AGHmfBe/4O/xtjk49nyJB4loaU+3AAuAKfazNg
XVWMTuAtmCOc49JhvMPd7672993689gQ94uvx+GtO2L9PQvyO9Tk0OqXj8CZfKK94FVhY6p4gkAp
cGeXjBy3QHc7omL5Aok04h203UskoeBzG8xRFJymfaUOPbiw2FPKZZr2frt0NnSyG7P3LiiNLkAH
mIZxoAeeYaVyXzCj8v3fhstcBlyAEb46uMoiGjYqBjmfL83m5yWuLZvADg1SzBR4jrCi7evbmNQV
2gtwbrlfJlxJcb5ZVMc1cMF8xKYChVzJteEK03Osyt6vb2ucw5JcPNeshtWHsHpyUYFhB5jyvH3T
q++DbQEy5aDQ7X5hfbfpdpRR5MRxR8bwRwwmsGzDidXZkVd/cM/2dOkHoyiBJWK8NEoUVNRKbwwH
SswrYDFZHuSLgvPn/2c3pAiF6Ph8rcpJeoZNLMto5BTaeBf7sPMJ2HTOBdDd36UwQKuQvmio0O43
b4Q0Vk4KwFaCoDKQtFW50HIPOgvpEUX0klHpI4hprprYCn2G5z0UUnR9iQenHIrp9IJCR54xthli
nW8YIfKsFMFHpRCi30nt9H/zKBoGjd/TGfMC5s9uI63jA5UDiXHNy3qhh4buUUoTee2rh/kLZr9t
pZH1qCcsZTmYUR/ljVrdPDmWGJ8KLhjC16tVxL0kljGKAU1xcCHPTc37i9EILL9U4bYHOQRiCrDf
mcJUVExeZhFXq1FXSjnNqUjFVNR0p5ZvkQexJNtVXVsQiozcvVmTe4kBtjL2G9jqjAE3ZU1Vm8ID
VVsyPZySlVPNQZounH4XQ0GQeAF2Jf3AhOt60BLDvJG3Af75aqWjZjEF39o7KOF4eQFvutzIEez2
8UekY+uj4lOy84jf+S26dSJVlwGjkLckJyxbA5PhMZlHkXklKSt+t3TMOk8SuekvPrQAlRngP3Zr
VudBCYzp68sb5k9LPzDEdJT9Ij1tCVJXsJ+6kC96Pm2OLBCONZ+2uQyLDfrurAmYJWxIWiw+ThbK
oCrKd1n6TlnHuzheGKT/wfwSA5h1bM2HxTZ9QdE2+mV6ymd1C5OQI1hAP55rGrYiGfssoXoo8cKg
cdPTzW5HpfYv04/AyP3cxlzmlw89yzDauAqS95cO/aB/5YenqKw1lCA0AOc5FBLhhlhV6P+Q5TEW
PwaN0VWK/pYVH8tlfTm89Pn+msdAYC0HUP/dQqh0nDTVl+lvvKlQGnpOs1N1yN8fLgLmJlg5xA3a
k5DUql8vfX8u/XplPnX1d+zoBbtKbqP4XpzbqJXeGLjztggtKjRId9OPmPBKUpgE6wax9SJhLlcX
r9jaCoTaJetJFkYcbs09z7v8yNTdqNfzCriGFUpFRB1kmIReNQZqMQvXjLf8G/q+Pwso24/oudP5
aXSmf/m3OWILaOuHIHepuC1SWClsKkxNXXf2hD2GuT9EfaWm4oaN06jhf/c+7tH66AqBSMac12f5
bPqOGrwhxpw7849A5umqN1VbcJdpCiZWL88QnvaE8h2S662bJnK8G++Na3nrHF/uugTPEnrzwMbv
aoss0YVsJt6MymMWwPZh5MWDc3jPEYWxKgU5UTRUeYCmKIymurdQH+w7I/asLnkBIOiC69z49OVi
lClCl3f6D9W+hpDObg0D4YHpvWPz/F3P0UxvogtYVIJL73sYpLuutY0zy0jNYA/42a0iQV4R9RVt
C2zevAki1Wz/Mp2FTAAsy+d2Sg8mDqCHrJ+1BHtREJsjjTF6fjUL11RdkR4HkFrM9ukWRdfqfCar
i0od4aXziwoMwzeptGlHdl9L2xybzacagVXkGCBcvvwEWh0LTaKYrCwwr2IUNgL6HTErR8pwf70D
YFxWrLcUExZ6rsakZPkqgA8nmJ4YnnCgZICA/9rouq4T+BWvFakA/27Jml8BLfSTeS/RUxf6ivwh
btY2cRDy+vsfsfXmzQXQL5e46B0gMpghVpu3QD50kX6l2wO8IIpcun8HDMavG0tPH/uM7Xyjez6X
iDVec0TBoCcq3A5OOSedzf76Am/yt+lkwMbMjuBXKKleIRvPgO93TZlhuRs9/EuCY3JPC82j4JgS
Syc+l2w+O0H+DeMamdQZJXJmQugpPb8Ov7x1we4TlOIl07nAVMuSjvtjYfO/94kdtEbMOUrpB9uO
c9vQvaDvqYTXl26ypmWfMn5J+JOQMnY5wWMew7nQIXFb/Rq3di9/pt02DB8UjNV4nYvxf2q/ThI0
iY0BdN+mmw9pt8I2RpX7dNBSRdA/KssyCpcW/ruJyerFkdwpShL/LdxXGjhdK1dRUWnBZWKJKAvJ
oGmw+XIjhtqr5ZnmNw9Bb0TD5q7+myyC4l54oFzvamkQ4EN+cIUN5/V8mk75zmCn5WTBs8hMsfeg
Br4qzmYIpO3Q5+3k1Fr9HOfds3DngIr5Lr4kBDho8lJhfbblZjscYHcp0FWzWr2IaBigESDe9LbP
aR+gCCvL3rH+LUQHsvEGDXPsir+UcORxrkOTrEhkbvAusYaImBN4ndzRA6j9M1h5h5j18uJu5NeU
ZzNm9FKrupcnMzhZSGrObCDKrAINL/XZtqp6JHeFaY2RzIxyguNapJfFX2cVqWlxSxokR7WMwck9
KmXZTFtpz5GKfj672LrVm/QUulCciQkpPtLp57/3tZdPaQkatWljI9tZTmJaRrU/sze/4ZVWr5uM
PRZpFmFTgzpE58CCwljR6czJo5KR5OCYAD9m0XrEx7YW8biet3ZruQMPF+4uTWUKeSwaM10qFgGA
hXX4dqwuXzaO6mDTHo+uGVi284BeQ060jdH6bQAqv8KkNV2/U1n1LWH1EG2EkEzT5SeAOW5u5Tij
wgwWOTsruVjUL3SIKKnKu8xpj8zUW6v9xjdmnKqHpMmkMeAkxoKhgbxop5UvghG2UUl+tb3Q0io0
5JZEGXAG/6poZkFpBXcWoMr8kIQLHKFaIG8WrZphFVaOmkj9Wv608yT2+yLxgQO1YBzI3VD6iskM
7qAjYRXR6/qNp7Rt9SiOQUnzdttUd/PkMKGXPrjxju2JdyuTCCvvMkxsb7fEZ/L2akejsIzod8dN
k4JVwuhguWZYpihXIXqv7PBdHiH0ypORTDwS/O3RCYIlJIG5wzZmSbb4tGGxVZsPO/CVmAgqbz9X
En7+qZiU+MM7jPrhizHdrECXsLpSGO00o0Q6/7xVE+S3NUD9pdeCYliEGHGQKR7/V3aUEnl8eVbs
2tDNnrrrdcOAhHLOL+cPQuzOLbjkXaI72e1mDxHlF8ADbe1E/Xnp+eoW7LoVhwTqScKjkBip1C79
n0Qvcuwk20AVcKKc3E3MdK18wllUi4wjtub5bnNzlhK7aVUTxIq/JCMi6jHgY4G6G7kykHStw+J2
WOWqijxclQD2WRlAInIFwyvHUh2f0KAtoHApNL3wMnHdZ9GhOiJjYvb9oz1NuZm7gVwpGJHbg+Rk
pxJ8CvHQzP+BFqsWeINkn/knv9KW3dFTZfn+1Mt6ZO5ERg55iyK1+tq97ZJ6b1Utnij+9p1Ou/nA
SDRluGcXItSivCt/y7/BBE4Brcwua0tArbz9+/RKQzTbkEtNG4bowVmMsEqnaQ2YXnk/0UIJvlLU
S/vz7HuZtjLEeOBghyCXYZgY0SWEn7FEjgNE1V1qccI5ZS1+5e1NKuc3VijIUEqZsWA4aIqeOJg8
ZqagpzqeF09QwvTz2W5VmqdgAekogDQoTqkY8hj0U/fVWxo6E/d5D4JzTXpc/HL2yqFyPmzEjA81
7WeIs6Ia65HuNiCRCmpzbFm+IabFNVHCPz1CJ3USJur7xSq3KCX/QlM60lQHrzZcZ9z5BpcINVxQ
jQN068e7OkOICmYHjlSTeOp/YReQStONY9T44ELGPCt/SnfFn0A+ZXBCE1+gh/4/BWm8efsg+uDm
D9rghim5eQuvgHPbA64WKMeqGrt+UiIW2oHA6RkJUs5/CUEydEm2UxLJdyDmKgs8wCZFI26IgZk2
zUuxWmMvHqrN6ZzHrfttXuXoso98AiXB9yzAd0E0RtkMrx61Kzxqt+AF8G3roZBOCwnlJr5oXJaa
JXnfyHpTedy/wNyglYcw+M5J6xJwEhuXnfuCYrpgpFCwBFdrGuP2nWjKWR4gbbB0Q1KI5OIxIJPf
6PGeNpt3heKlf6+XRGVmgqseL8e5Uh5iMhu9Cqt47YrQAZCdQji5H0b0Sl9GQnVh3EUHyUWFG2Go
Fz62vo167JvPXEGdopQfvihlNacR6jFyYj9RkxC4RHzLn49Nocn3I4bl8fovwD+OFk6LBVjpNtp8
evqmJ0dY0hJH/eMVYB/VGQi9XBrF1ETGnUvx+hynXbpmprnBT3obnuL0Z50FhYFKtaxyUxTcMVca
3c89R5e/9jq7KTs6b5aTbmHYYVYTbJJURumIZ0ctWYEKCrxEywi5qeTXCkELZWSBKOV1BBIH1e8h
/a/0m2ya7fbu3TP2kBtuP3OtohNhKNFp7THE611SB/ygKPSszuLf66WxSKARSO2xbPyVA1xDY2Jn
9By7CSiNhX8kh6XmXjMyU6SpIH3WmzdhxT2eu5+zUpYqN2TGYwCr1ZC7F6IHx84lZq4LvLLrFGWS
sMjKfddShP9pHGC5vUKWO5Mw8IfBnWMobFfrtBr+UaWkd7PFDXpwCBeMC2ZLnhDxsjgg2b0fAvk2
xYK7R2ppycgu+fw4DmjZFUEnZ/SltFpikuKhxsv1POFeWAfWYoX9XXUOIp0uD7hhaYyCEl6gXGZn
Eqmc0VMV0c1HfdFxuMY0U/nEVQY3Ib5A1q+S5as0CGDJK2jlGB3yf2CYMCxsqgzZQu4sI9M+T6J7
IilunIC+wJs7VLBC2NOQzlFl0MJrpXZWzSICV216h/XyB+j4bEpWGyZOQu3P4oK/NT9qJlaPH7ZN
VvHBA8qhHVylZYIOwmOhx3b2ZjK9I7nE5j1DHjsb/Dd7LkldDEsao7lr76hb2FxAxYdMmpBP1mph
kEVtg3kGg+9VKk5+xUP3JuM+OjhAxifi8RP8qBLAeVd7eDCsyP5ZETP6Rgs73NKKPcM2+QMj2jnf
sO4a3ESsxB9qmz7lDUvxEM2H+spJ3GqzC1jzvtjp5k50qEIBKT8JkCfXR6Ww6DyYtgYC0RVNho52
qxCTpRLG9Gmpb5+wKmYycNNSA0COyMdhwirERnqNTyMAZ2Vca7PKFImvXuugapymi6A3wmxkJwRY
sp8bZCgmVe8Tqbj3KZ4z+MMF0BMSjXGXh9z7WXJ/ftkNqHT36i68JxWl6b1vBsCPJ5oYgkRTSc2l
0/HRNLkfMLtiDRrkmeGQX6z0hcQTg5LjqtdRfG7IouVgd8rMIpK9VIaxNqt9Hxht+gBq/iscUBO+
RiVWRD8LBjnBnxnVxTiI5nLdiocgx6CphGXR2fvhftPanmMxqOJgBUWyvE0fzaY41IJz0Myndgg3
1oVVDLwdGvoIXhAhCzubTRNcFN5EDtWq3rPWy4gF4P1+gpkvBvR44PfxQgc9xuELvApeJ3C1XRNl
XZ8EMa2P85wCBLCt2PxQviayDBbqWxybgetY3ccgWylamAt7HNopKIu1TYqh1dle/6nAvksW/fLa
P2vbHTrDklsmRdcgfQcswHS17uIG8wbU27rCdvn0/JvYSFsq3sFDCauGxJqvDkUL/0QZiC9OhFCW
VpUc+mA/Kf6AnNvHEBZt4pKz2ONskpYHMORithg38sELtESJQHIHDQw8FldqD7OAKfEfxNMY/qqF
ZKLU3UxaZHr+l5OCKXUxStTvxvQfsvX1Y/QnWQRsstW4IVRsK0Zgwryg3ctDGcTXNKo3T9nWaWFb
0g2c0XazgWCEG+IQUIGQ+C8aXlLDjNDCX6dpRaqmP0PFztgdujAi7btl61yHzr4ZgDubRZcfAnaf
amv5DBI4IcyXyocWICdoWTXgilPZ5Ah2VRyvck2mu5+fMNMb1RCUzm9Z+0v3qV49G5HN6wWJd4Qx
JPzKPcf2KH1ksi3Z2S/niw8Avi6chtb/qccX+7UPseuCHkyeaBsUCSNcCk0u1dDhYP9dJ0nhsHMv
mCC45qsSU1KZ9d5GvvcrgECKEdoOrTxgPrEHPbTNsBCkdhOT7LcluJg3honT3R5doAa0NeCtWUCp
CQxpoxGc8shsrYQb5i3sQ8mbJCb2Hhxt61a7lvDwagh6vXoDKn9J14aP5j2SKnjzvUnXUXLFlVAt
HFFR+pDx2bhoElIV6qaSESTSRDlnHj6pRFLFsLEZEcGw6SCOp4D/gZss0sCRl6AUXsmRK87UvKx4
zUyZyHHaEZxdu6DmHLAVL84lfSmgij95WAQqvLiPLIr1e+qaRLvFvkLw7eeQzDskkQyDSmxD2ZqG
j5seZkTO3gkWbXg7Iv0zN3vC4wWjPq+HBBh1caYwvUfSpH0EX7esZLVjK+YfU5BTMKE6Or6BSccQ
EMpdWAWv+zuG+Jtq+RzNCCRiQI56jE0pkOZxd8E9bIUvl/8HR3jk7oyWqRTs4L3LngaRcJUtIxr9
cguDdvScvEdNvr0u5C40QUO9FOBFZaGqFYZQtj6U5OhvltsNfoT8kVCgq7CHtRbuhrVnjSOWvJLl
BBioddvnG5Xe7EAbndUiVbyTEu0FIOib7RLrV/CiOIdb4i3qYPdGGJ/TZnARWVXFZ/6AcxnrbrBc
bicFcUBZ6rSvft+vZYCRBNKSHI6BWj5H/y4Byt6FHPhh5Csf7aT+8NBgHvyz4xPPqGDswN+7q4cL
cU9OH6yx9liYlw+aiSObivmbIur1LpCFMIyOFmvle83JRVzrVbX3rXWyT7kxislhUEU8q5iCVEg+
xn5ocaMJ+AH2FX/ZQSA6rTHxG4TybWis8m3JgyG2dcWiV39JKRZHMeecr+746HB77+CM/5B+uabt
nFywxg5MHoxY182Fzl/9xXufgf+gUmvqwkQqsForoZiytm7G9QJ1sh7ZF0oj8VuJdAbT/pxl/prG
qy6QK72IbpbKS5d0pqvn5pp2vxd7wvM5XIGtad0ZxthOYrCvY7rmhpn0F5FgHXqV1qKMPxOBDwpF
UrnGbxxCDCkax83JbdhfMwp9b/c/3Z8S+mkPx1DIfnnHzm7TJP9C9vA4uJ3nLPvMngdRZZtPEKFy
9sNsIzOSPc/AuBkDm+abz1PNUQshVeEs6Sj2B3irv9ZUS/k8teI3CjW1MSy1T21Vm3nDVrsgUXdy
6fg8eqGN9bU0UX2lny6NGXW/HHz+BoXahUI6e56INBYtP7fkpYBF4Hw+eR5RRz+6ECtxhbrf3/U/
i6ppHRVRlNwFTaIovDpgNv071nLVfv9cUK6qTbhIf8xqNKOgXlXu6prpfF8leBlnsgsjEqm53KLR
tu9VE+6gf3/oKx4YxjXhaWoKcLj/XgvgSXs5H6X9Bv9QffhNe8Wtg1SWD8WwCWnoMLIdzV1W5WZF
RbfRb3fupVGi6rT/On6MeM1ROwiZdkN3qHWjAHDM3SSV2fF6arf6PoHurtCXLyEeKKwPnF1NUYX+
hwrifThYgC1Oo/SxQh/JcfTJ9lEkNhEQE6FeXMBbluDrZAmWRz4khjx9afq82aPIdJO7q6X+/j0m
cNhuWVkuLzogeubWWMco1hgksLJmz7gqxUSQblb4Jvdtji32kDKiWZCXC6VB11Ff6PHlXtLfNwoi
NQKufv3U5R5rpcEwi/mt56FC6Wi3kT5L8/K5DjQEkex75Dd3qaDog5f0QM1RSpkKiMbKuY+27fd3
0rbQEdCHWA36rzUmXgVKhl81cZ60lRcsNacQ9y+5qyPReP+G4Bag3EPiWT/bkN4IWCqNRYJb7jGh
MzsF5Zmb+K1ooUvKLJ3Ku77izAJk5WwfC0t17m/Etb4Po+W480dciCrqAuGOVFGc+LYpqng+yJ5t
vXaa6QG3od/PM+bIK6s+W6fFeL1q0zGNyf/NCy1+ifhXQ6hnUFksyv1y+Cb9OTTxM9HhhNIXfDoS
z/kKtlKxgLRcqtGINRDeXjXs18nTxyjk0/TI8/z9QRhnpRfOs0CIniD6FsgPRgCwcgWvOOQnsq68
20xuZIFn35+C8KLTLJfgLJsuRNEC3XK1FYPAC8clvA9Z1D5vyD1QUSj+N818WTxX0AvaLDVnVMnm
/BGBG/j3UjhmjzPD/5y5XtuzWa3n7+fE3TvhpwiAWZN82jdw8FVflxqT4LzWJT4XZRPD9n/rTFI6
/Ztf4+Ng+kUAK+PPkZRuMOoj9rSja3FzayQH3saN1XwVa9Sfu39sZ6FNmx41Wj7FWG+1cNRM9dxM
wHj1cUZIb9tIkrWUNI1Nck+rjtcJaCuls0GArxUFX7e68bIjei8HdytQsiCqOahZ3iEvczFPbrcg
UTQzFuuuE1zFYB7s/hK8uxubrIzrF60VMfDqLz+Tiv2inklTf6KrvICrBf6KEk2XIOb2ivfW8Yqj
KOPfbplTjr22ocI8oE9xXRiCsWc7VjVCq6A1cj8ZvZ6rW9uQr1x2a2OnCA31m5LAF80zNzzwRh7n
1BYpu8eO5tUtGk6XhHSuhT9EGyugsTfHyhEast3Z5bBd22moDnz3GUlpZDlTt4mrpKaKepWWzs9t
MPZBFbT6sfzszBajx/fu9IG15ACI1UJkVArYa2z3LbqqqM0+1uJ8UWLbvGMDVWw8qXhjiKtAAZfW
3NGf5AfwTumdUWFvciDmGnjdM8Mmn/l0EeK7U6xhnvFpqe8ZGoaE49DCdVv1hlG7zexMRHBkCpgp
dpgXF0M71Qv99pNiAlOG/1u96wXF/A95j7zU6Sor4KKczOVTeHn2YDnu7d0e1f/8w5tC4tUJsbcB
P7MFsfZVOUZ6VFQbJt0O59TSCfrkDwNsBSBNlgNbSzodJDL4ZlgOYiQqqhTFdLzpEs+0xA1ElNwy
6Cm+E3RmRmvPxyB83cQq9DN0I51IRXoxylfFdBwxjToCPAy25JyrFF+QEzRJIIK8Lr+DpGHAQgnR
fY/AryA/UVMiaPa7TnZShHNX9s4cwkegcXXEru0ByKtAsBfaWD11wUKJQ0ryoSpL/VFHV85fKjfD
1JmFrd2ZiFOcrICeOJRyQCX+rsAnpr6rakakdTkjWoAzGZsgNQFzJlaq7aDf1o0jOcINPPYSZKS1
mdyo6j6q6hCVS8iWPGuBDbXrHv8ycekuXrmo9S6uyf1UIDVYOMLqFA0DL1Yro1NgmZVdK042fS2t
fufjP2Cox6VAOcU9mXPnLfFIsJcRl5PZLSJgQ5+yiGTgY96bvEG8nst8z9zai2Q+rCA3+XkhvVAk
MHA+/gYKbyC2UWtLxjOng1tNqipEqtNHNAsip8Iat2WbdJxdUgMoQcIt/l4W7gdxwRu26gk7DPs2
JKqLba6pW0+EH2tCJCS3sBylRqt32OOtf2SBKt1itA93LMGj4yQVrgEgtUjQn5Gz+MoDZDkbUihJ
vkXjsLWvV03liCJz/idtoHJVB4t09s/zihDr30u0yN+w3J3mcUuzJJP63JfgDGg5fQcFAnUN/FRb
XojdrLiH2TbxAf3uUIMon2LyYtBzNGqhpilbjmoNfEX88Ay80bDaZpnmeUt0+JBchYwytqTqHiw2
KC5oE6VT9Pn+WEQmv/5Kc9iXAhcRzxT8BzirpBzJVOe8+yJ69iZOuITF8OrJzejjmHKlZarP5fiB
bYekengo75fUz3L/l06K3MtScIkoKJl4iDK1l6EeRN6KRQcQv3Dzv58mknl2AplFrRS5hCsEdOeB
GGHWT1MOoImZ24TXo6kabhoT4zZ9uebuCwkMYFVAicYeLiySl32YIWJgMLGRS4rPDBtKSVmhtMtY
53CpLnVimF4KfCsTB17BS3YjGC048k5Me13aOp+qEHuUA/+0w6JjP2j46ZJ8y4w7rm5ABbx6F3qZ
R1vPGwAK1H3l4yu+bBHQSZheUwHFlYxw8aKblyCgM1LpWxd4Si6j2TCZ04AMb7jzS4wtbncw0Wq2
+9rwdKHHH0eiTRlAzDxZPGCd1ms/8puOE9wMBtwQRQG6UINm3EAqCzUAdF/c6hQ/s0a9VsJx2709
pqW/axK/uk54t+9P+bimKLXNn/WWnjBD5cjHIaEn7A5tKmyPSBZcF9ePdsKpzAYAohKfI3ImC4d6
0mhMU1tLo4BZpqNy7SdlcnG7jTmgm7ebgD/GAiNkamrohwiQkThmJhenG4OpO1iiw/gAQRp+HLPx
CUt54eT3LaAAFlIoBUN8pMlqP6Xr333FNUiD55SItccN5FTMhNw3GOHjs/aGPeVjtHQRzS3c/GFs
ocKvrHCJJANJu6ydC4YcjDEOEBfI38WPTUOxi/9tQD5O6qJ9l/0ohpK0tKAXPnMo/B8ui9sAUf5n
i9/tv8pGv3K+0UFSQJTl/+8eZnKHYi+YaeakLtDHt1T0ieyCVwEZpWHJaO1NX7eDj6g5AhNHumsC
Reqh2iu5QIP833CWYKx5/09XILvmCNxOpATkpx18s1Ol4lGUGu5f11xCII5T9EiT7BDnNyGSbMvb
b0SXbNHmxVpAGkcQU7qeEC7KUTHk8vKcxAZueaRzxbRH6AE0XTQhAEXtFtEtZLCAV2Hhml3MIdj2
tJxYBzeKZr65/koxgKj7S125W+ZyfLgx5/Lf7+H2VUMHod0GFXrbEBIZc30bmzeiJgirtCf8sKRs
qR7DQbJQ53Er3BVfKPYpMYnLcoXxOYhIs9dJ3ZH2xhaIEE1NSxZGVWbT7wCunSn3okMaqRwxU7fh
2jghQR8nQN+prhHmsY4SCe2pbjmdFkp+cVmrek0JsdxaIMYHqnHcSsdrBnFp0cdhLJDlmIkIVr0N
wIO6bYuAzT5Wsr3LWKuWkhP2Nbdnc5vRMm+M2aE4qlaKjsvcXmDfDXuLf7KimE+2zm3qngOCvOES
UHcAU8N5BAd/wib+esyoT3tMgaPyvl76a1iXOSC5VEMHee9BsFyw7jCLFeuDjdVeTrUHDerLp7l6
m5Aoxkzlh285Hr6/TNYjr5Kw3ktGfl2vE5BggNwtIf9nN9WXM7ud8PfIGJ2Ra5KxN2dwsXu9dJVe
Zxp3LC6I1QX+cnGy4uhOVO8npKrSUMOj3nYI3DNX8T6rLBxyzfDe8kYAxIqkA1jvYXNU7uMoY9jo
vamLWTtrMKAAS8wb3cHeyTq+ez2RUN2OeH3A2kx5or0rlX5yRX0Ab/PyxI2qCl2C4FHpTPUujE95
2VAogAkyPy9qjDwqY2aFudvblFYnGvECkVQU9rCK+PfQ75x5TiKQBbC1wBVkWvrtxB948TRMPVuU
ZSINo9hWnTdB8uIPYLIkqSsAx8Yt8EKlK3Cp1WBcydeG+7ramPrBgqNIITBasRA2nOQ8Q2abaEjp
nl24QuY7KPSaM2Ds8etRZ55FtKQYC4Po9zopcjwCwifUzhQHQ2wkAWQc3p3D8aJSx/25dfJvEZZJ
YK6WLXJg6TOAyprg73jQaGIplwnE0R5mnUxTktnWckkXGRmTlCHNSDCNcTEFVH3eq6pXQpKr6K4M
Z/nDFjwfXIa8ZMxEvhMWbnjuziYoutDxHneItbM1yvI4b0uSBfddYwfUzJdQHGyBb7mVpge98ew9
uYPnQlEkJZWBFL9XwrYR6qkeQux6CW9Ybs+1rXIriKjrT5dtXAezCPYnHlZxCISo2PCtlZTXjnIz
6wmlIA8mSflB6HKsIINj2JR+EjgKYDELLEEbNe0ymjdf9XbSt7LgcV7YQBpsl0sjo96xxvLhSND3
3Nrc9CZJU1TB4OUnmDhfDl8Vd3LcTZzZNjaVPZcxqeKVdpofzQKlYw6OSdX9FY8acy5xn5IUx5dl
aKRTiKauySBL+waJujWZSJrfvdTZ0UVLICOc9fBebueMffgYDr9Ac8JqonF/HDPTGZvN/y93zRWx
o2zzdugHd5szXGObYkiUUlude5SkQQ+PWeN3AIU4A10ZBFfCS6xqEgO5HMj1eEK6ELlx08oNN+c/
kxjfP+/BLg0x/9J/EDADMRudDWrjX6LAHCnUO2/Vnis0TJ9/fKolgbKTJ5/0YcKBfCWP0aHmimsL
nNBYEdZid3Rg8bTBkwiBe5Pp+bt/oS667bQeyWo/FnNii6cVbhWhGaNKTCIsXajKuJFj946u5c9J
KVmCmmNi3+KEi/h+9CPPc3SdRAH4RZBpoKE0g5mS6KISaJ5gvN/RwhEIiUQSTyhPuFV5BkuiwLMu
qQcKh2Z9mZR93TnlGf1h8w/jFgPv9QkGxyA3LcqV9LPGBaRgAgzy1z9a2ffVIdHpU+x8Qz38c7Dv
cirX9lUpKFqlYfwh8Acy3ll8nUaYgh4+WnamwM2r+11m2aCJ4cXP++2+s6yN0zS3HHHyUpyqp6uG
+qF2OwVSMYB6DtwLqWSS6vsj9EpDklGhX4pzWorB8EdGAkePbj57X8sajmtvT6CGr253WKZ5Gk+f
bX4mus+cHLCXzB5wjjb+PuklzZeMSjUPPMy3t8S7DUso1ZKhyRlZzoTBlYkhmljBj4819s3vMqHo
SorxmFixyTnqKMyidZzdj8Bm7v7mYBf3xO4y/QRxhSw0CRmGTi03clBi2aK0EYge/wI/1DXYh3YL
Pp/fat/1S9MOJCNm8A1VcMqVAY/eJN/H3QgcdJidTFzUiGbCzZPrqPLfjzxCibdGwtItrGqoyHUI
MR8S7kwQHl/xJaFZIGWmdcC5GgPzVF11ixFN+QYZ/DnqI0hMbtFb69A4C6cDy3CdyNg5tBQ+CJQR
QtA2Hix48MeMRN52F9Kws+JbH8s9BnDfR3GUK6aB/E0DgwFWBP3V8xy7zvVqN+xyAGb+eKHRBXv9
Mb9gchwXIHMBKsILh/NpYluqdgivNT2Uq8zED61JKvS27fRi0wEArixai+JdDDD/bsmMYn2or2S6
GKYVV0oladaLcZqihk2ibKSVCVGYsCSG6j/sHgXgcq6SxtmFtijyny+zzgRq84AW2467Z4jPreB2
Dxjb1g4RXzVVeJl48Jul+3li8wqUkAHHk30mmFUVVrIdQRRrA4CcfCty88LxLraHlUO/VBZQTREY
6dVMAprmoJTsWqJKYiDZMGM/gSfHuIS4g0msRKGu+2JLRZNg1aWta3AcBLcfBMx3TkEO4TZCmxI0
IGJ0C/VQPOCezEOPcQhR2RP4OOZxyxgsQfvw8iIofHTnidC05M63bO0k2zhPQ4JN4cgqjV/5ldMo
8D/KWLMqXqD1Bsnzh3NfwUx/b09SkDursCq3TbEyKAC9uYdlv/owNZWlEVGbMdsKuqCAnAdurnga
Bnh11sHsuiTi77LckPEGbp/vcQWwaKxkCnHQp1CZs0vOT9WzPvLMJHmKrmldhx+4hgLb1t2TJGla
F1ivxmaUdyvB8VWEC1fVW4Lh1XBU33Yl3Aigg5da7cL62gvflpAo/YGNPZPl9BxATkuWkbHcDYi+
fZGD94zSd2u4/L+y3IY+LF/+LM+Z7G4SlogLRIPUS2KHABrB7FjI3nVCbOzD4rHY6vCg/YFj5uDw
qjggjnwwLebejcvf/Cz9HXfcR5zYuvoR7TI7XaFJj3C675KHeIMz5tSGuB+rt/KzHSpJtqdoHxht
XcJ2JWUWxukNRxRmiEogrSiu+03za++qKOZzhsNTbF0vvOavQued/XvWe5uRsSbXo2PZmQUp5WQb
S6tAS61ji1ph7EUuj9Xir4OVeA8b4Ks9xbvGt0ulpCU51/uI9yGmluVf2mPwFmoBoaqsv4W3aaOT
8tWKGwwWcKAWXRAmYcQs9B5/L6Vu2i3jayiohaqRfFszWqiO0yzYsrTSCEBKdZB2X28S5ks5pr50
d+/Vm78P9upXoRj1dJaulMBkheHTAlY4m42iP1VLi/jgYALQ6OnGH7pwM+3Acu+1VL02YkCMiAlW
HlkmjgCVwloFSlMyAavVfMd7Tw9cFXjLaFLIy0NvdAhlpoeda9SV7CmZLzqwiVNCFhFrv6pKbGOL
f9Ci/vssZ6N8a3TgCG9bj6nkD7u8sihSc64UkA6ByybVbng25b/QfK/sxOEKGgFdkwoo6Vmjmf43
Aj2HCVEkTfEZJCrGV7dOWPqjs06WoNBEHJHVKfI+L4/HTVRtDamv2o6GiH3MyXqYBUUNhxjQfsPY
TCALkLJyjC9BcQA88EsjEHl1TVh3SUo5btN5WSrdfPiHpUZKQZMTOD7oWAD7U0JZ0TZbbj3ihZT7
0/P9v7GhbGgoiw8PEzZbtmW+iFA2MB2ihxuAfLaZNBnPi0geT7EpfF59lnPAu9c9XsJDyWVG03oI
bfmMYOtYz7tAtCji+fXqBCQGECZmqtH+O1GROyUf9GY41ZKekXugLY1LagARsMPX8LEjaHYnPzil
iXiBm1DgJTrlCP1elhHR5xDkEBLGlyylY2pjUIuU+abS/B+WNv9mYp1CaJrKKUp7R02T3wttbWJ2
arizeXWpdUP8h3LH2pgdoAnRMlx8AOIXynhxTr23GNOcfdW86Va1nxG3fba5nEkXcRX/Z3gJiw0a
6dYj1fo8UyQUH5EF1PAS5zeRC55KeLMIPqT4Hp6eEMYBwjuj6gGfE413yAVoJCLotDBmEyJGD4LU
UUlnsIUTsewg28HHTKTPOqdy4kgKf0Z2qNveRH12mCKyX9NToNvDAxFkhja9d0CygFCHb+Oz+SkN
TRaeoT1wvHuHtsjQ2uY0pWTP5/mzY/IIUpjw27XLAzvf3i38PgKDmNJMq6u+g9+oRKup9m0tB02F
smcAqFRPWovaeWy6XNm6Y1hsmehPd0JtgtXKT/5dREJPbg1GE8XVErMMlF4ECtKI0jpxdvzyOiU2
FNJ4s8zYSU1MjQ0Q6p8iaJeVp4eTfhzQvSi1O5yIe/NDqxJVjCaaIf7u5jd1a4wA5KpzLaZegPzX
lmd2uC5vveDy4UK2nTraRA9THtQd6q6x3+5Ft8GTi+5fFlTas3Bb5x8st4g0llEjcGFXgqSaW3X8
qpURS6ubXg7hTDNT1+2kQ988+nTucmbexSYiC6RAwOKv3YOrNzomWr2UtDZj7v9pTv/G/2YmtyUW
wlG/CCrewdk1VuCJJjmQYj88bmt7nbVjRAUI7MfagO2JMSLzs8TJBJkh5XApCrrpaJVecsj8Ns0d
tK9LAP0Wzy/layDsNJ+Nzr/rg28WSKYywRkd1YImQrcnfbouldDcFiCd3mECUU2FP45HJgfApbYm
wKSeSg+OoKucWeYSGmqb3ytEZ6UNqJ2GfkraJfeGquKZeQoa+W5hxBPWgx6zRZPgC4d2/wRiBRDt
iwhVUEC6AF9D/UvFtxNIZD38JkgoNo9HKBRO6LfIchEdGqaGgOboE66zXBIUgh/VL+y83xo94OqO
HH91JqP/WVFORiwbMbhfE76A8BjsCeyiIm5c0rYSjPPGl7FGpv9Q313H2jioB+zSgR16adtqDGgY
5becsBx4qFJOExESR+Z6+3sYHihM//uhwt8OKZhCYE4fFOx/kAnl4BLN+Mzt9G5KbUdfrS3ooZ/o
MT3iVeWEiHqipc5S2xa3rW61Qd0zvo19j2uSnPAgZySY42L2Mnb5bRocjn+ResocWTySuLbe5l2e
mKvsk+l7uq5BGFO/f/vbSn3LMsjM+w6kpfiqWgsuLIHGpobSNAXlHcze2aW3Z8wU4e4XaoQEUlS/
rHO/PxpiysMGmGVBucitEU9cwvVwaPuw+B2JWJE7bLBQsR8ztI0X8y2MRA+I86dWWdhA2cDYMpSq
r+SDdtFFjAoEs3m8ClJ9FgM/BeaW1P3rjn+K1CPGfeKzYMe31qjkN0oxE/aaSTjTeGBANMoENZ4G
Dj/9SnpKmYNDSfLiFF8yblOU1DchqXlDfy+T2r049usW14quMOUIdWIcVkVDlcb6xWSgCjWFosLG
rhFrZoa2OmYQhyBVmfjkHzTw6bwI8haTySo5ItuwPJP3ZupgTbKe5k75dqIf56Y7x1firLWE376P
c1nixWOQo+lbutf8leqq3TSuHCu+Pfnt7BUKfHBTQMUBLtKNQXB19T84H2IPxbLzI5VbMK7dKLnT
OchDshOTu6Wa1HXdyM2a5ahjH9RXwdiUYDb8kA6gb2cQOuVEIlT1azuHzJDz7giNule0hcJCWFaS
wKpNBe4d1LTT8oOf5ztQYv5KLIPi+QmQ1ERdQ5eN+99QK/uNcqcs5fXQfQfvyLOGDRNbvE4z0HcI
f+tD/sE63/7qmmjsunFAzOpe0Fo4Iqhaz8MRQkGh9mUALrZYfRiM0Tg6o7RUWYfk4yVn1OXAQSoS
CWoQGRT7w0Fvr5Uhqzyh/pBJAwJdqLiKfLdgC4nRzq5+//waHHGOnw9eMP9Ai0bnQhnVm9H3c5IT
XXnk4hu9XGEhm2Cj8UHx/LKoFWTrffjpjkGaI4VMq9YVhSutNFiblVvxwV3NPWMdxTmo6E3y8CU1
qVhnIp2AXddaJ+tA53QUQvc4zjhfmLtIgWyODVoN+UOYyCul2Nqbu8hG//r8thwM3hr/AS42yuAt
wgor7H1hb/d5kWUU9gfXemAnhK5/RF96GvpsjEMYJMdf7CxgKFqU8oiy5HiyYAbw3igPpfX2246B
xjO5sCX0rY4kEGJbph483yxLIumZYcPP66ttljtHH8HhHUNg7NzKAdRaY7UE0YDdiLuSNRquZnH7
3gaadw10Q3MYFLVDIVMsLlcvepoaSuJp98OjIR/b0ku76sQPC9wgZNaGU6YRPCSVb1ytin4FGckV
Esn9j9Cth51jDqXubbbXc9KHxtthTzuzxwtguisoGEmXc4oyzh2Kccgwv5CMWoCCrYSa0A38G6Oa
jKnlVFVzPtMOf601ca/SABS/tS60kMCwrEDrf5uElcK4iYu9dXruvihckQ1EaID2TSm8z63QxmP3
Fw+3Jz8Jyrukpu0+eWljw6sbnX37ZZRT4GOlyhxXabVNTcoZ0QO89A8kmGhbceJ6/Fe41MSivtrW
erwVdbonBliNz/7lEmtBjuQ879fQECYnwa7soi2FE8cCvuA12jpHTqLjxZ1UWQVNedWoJKiRrtqN
JCDWlm+H3YQFesEQag0umihBe7KOUHUazlzIQSWr2eIx67xAYS25zB6ztReQAIbfOXNPeueRX5DC
sIkLhFAEQWwUvQ3Lv+mGGLjlyl9AfRsmiaPfF4A+bM0Uiw7kIZW8UC/6+ImtUuHr6hmj7EjOFAL1
zx/V0Yn2MEH+4vWb5Pd0eReu7CPLH1Lzr6+Rqp5C6Eq0p6PNLAsUEqwIAoVBtL43dzKMYEY1teGa
BPU41w9w2LYzf/uFZ0O7UaEmMuaIfzjjRRxkkrcpy4Vsy3WFV/0h9J5FpMtXCQHKh0cp2Mwd9eLS
YnugfbfJ8A/2ZlcdFPYY+bHzFM16Cr57RRLr89vH9lVU+GBpkRtqDc2eMZ+u5kRKK4AvdaiQ7Oip
//6MmgCfeTRVKaN42e8J27a3ASjH1bhBx2c23ncXll3PNRPePS8LUENKLKz4IUKbQom1uk7MLu/Q
V/8qbeZP2jSZtvILUuTVrQ4NVrFL4ulZM4/BvGfG38T2Y/ZyikmpO7gM5X8VF8DZQeX/RWyA3jdN
CUHmNDnBTs8AfL93udyCUCHkgNYuJShAXdM+BkkN6bK4yyJE8ngr6vrXLifyDe2FAfkriPURoZ29
vAoe7xm0dsOMiNLHVEixQBluBONF6xij6ZUCfIE40FR9Im56pgj3FzCFmsHAHIljChk+qVAxc17M
P9ft/EGfIn6uZa5rVyKAyLrLtEwXIOsBCaYPfgHiXN1r48iY9AiZAU7gdZiRSpYgFlgsXVUINjYV
iiaDxYHWKu0p2qyEKzXMq6rfMHeb2UYQrJd9yuMIuvNtFVehUqGv23hKQNd1C47APEnJzFQn+E3c
RkwA0BalbQR6Rrd5BWPApWYrXIMOOsJ6LUML1KtPfr4HNfNOEsn8yKcDHQQRxmWee17Ny6d2Z/mt
8HvXIwWZ/LfKlR44kE1Hc2XMZ1ov0tbySq0pvfqmMEA8T063+JG/3TPAUC95sLHL0UO44gp+0v1h
mSkKzF2AJlAbXiNLlIazIhjF6PoqCUXrNmxCB1w8x+iedZmi6lk4egFr5lmLyIwTRCGltitMpCpE
AAlUClIhHyGgAaEQYyWFxSnojhXtEFcsJIPnc0QTOTwsNktO9VqIEiBMV4l3g77SYJ6eyIQnIcIl
5ofLiH9XqzsBStBegh/eP0zlPe1jiS2a9AuFCp/TP2hgGQ1X4vA//2O6qDbGLYndmpxZNKgUe4My
uwkCwSWZvyyOflNv0qKdamF9WJbDEYumCcf/G/T3/rPX7YJAadHz2Q+1rT2kqrhEL1Y6Qw7sSl+4
oc8HrpO8OgffpvyUzDgEgcXQTQ2UNzQ+tK/TydqqcJVGRnsztdWYufqMIeHShiJt/yfOKvUfw/ia
76Dv0g94iG29GRCXh6f71+Dof+itCmJR4ja3bAJYtbtNLVcDM+lba3jAmzdtULkhkusQPHJQKy7X
xm3sz3VnsuuHul++QFnuw+6bEeK703KIouqtqbPYZiJ8LXM7KtoUC1Zk55ViE5kTPB8p07uQR/XL
/0a1B9A2MVpyx504gXoTPnqXX3k2In8h8sJ422ZrEsb37e6sjZzaf6fcgDPUKWU8C/LZM42g0CXP
FuA/MYmnE5grSlOH0a3kMxOv9KtqRoy3eHqTutqfSlOKjgNIDCkA6dYwaqhPHKXW3huvr1UZZzIw
xtzjduZkyWIk6VAmW/PBrTUktS6Qf0c+CZByX3vRd1TJBpIQI62+d7DNO51EAsdFQDQOG3mpZH/z
PmxKob0EbSz+K9zHbMqGJLApNDCbUcUX6CAgj5rUxUuME8tA/XSLDkHkTTxZbeWG0beqFRhubhZ0
Lt7YVE09RFXc6U5HLuQm2NJsxea0okPQtpxuCQArx41MGdUtrkCIQrdpePWR0ZIpUMigOWkm0Fx9
wxdu214r8Nr4P7KkHZEVsRWQ+2nR4lNAtpynjAxzpGJyIArHUJ9WpPyDS9KKIjbLcXHtsnwnS/TM
+2dMI37cMsoYOsEmhUxBSBQoQvUe+n+jYCdoehgg2irQ8F7+Ifs2w0m2TOGY3DIRyUC9mVQgpqEI
WTTc8gFKOMcbXcGA+lm2GR/uAU+9UFI/oBDStNewCzFCo/pv/R507eYSsWmbAmoVjdEfdPgKE4Mg
LT6iKVowKEjAuTgwaTL8sAkYpU4p1piHCJEdOB7jQccFpPk9vN1a0kdpHLnd1qXu/6lFjBRwQbF4
DDOSq6FSS4WM9vTPiLQ5j8TLkxYoJwrCWKJu6fzHIY8lqllClzShS2X93qDD2NP0qPD193e49W1m
NFkz98rbFaawzlmj55G4ETzJJzynJ6l4qimCx7D++JX/75NndSLmnZz6Q5jQeGSEdINNv7qJcVz0
Mi2a2fYJKJ8KaC8rE5/7ilD5injXkbCfrDWYvLex2QW8E3rkUV50DaqCb4nhAzzfjnHRLgWn+pGs
9FDzNFdl2gzOfhhWhDCAu2gli1VJgIhhCg1RsGUt/rumzAMlQjXf4CeuuoFc3m5bC+6UqrigzySY
MkA5k4ruQBLXsbt2cALzI05YPdEjV69KRNxgeQjzFe787ynBbtrY9Cb8k5VCd+ryEjvDopz0b6xY
tC97nx5HI7eCpZAsPXl4ng3fYmOwGCpnT8ls2xCycSBb5d0ln9h4Hi3KkDL3MVqZr8JfEHzQ8yiQ
YV82RPmj9baT+emQ6dLMHy8o8qq9vgjIxk6Y5Sgx6S02Qt5jDP2yImu4hIEHLF3W3F/2i0DkDZaw
xUwHI57iJZr6OIsxYc0XdajuU/0PZ8SMX4Hg0hy0pnKWNflc4s9Mjyh8+W5NSJ8Ll8KzfedxomqO
GLEhfTt4KcOAvIwx1TPq6DufXe5EuUql7HfNpBLGLUhcxL5UzTnes5/JKRVL2GKXDuc+yHMJnRNI
gc+Qt5qoDaXLWcjkK0heh6QRV2pvkSMOXNRbrQtYQrT6OUHOX7BRZqd2Yw3b6b7cUPS3X5VHqVjh
7gHT3Q2VoJAr55JV8SFcsvksUG7Asjb7Lk9C0q/g8aEkAtquw+KnhP3mYCqoRZq+ZN62+U7XFF98
VM7IJymmeeU1CVWg2y8x7xg9vPlvn0WELqDYDM1BXdU3/9e+WrfRrYs1AOslKmDGz2qq6mzJ3c3Y
j0yWW4KP9Idwi8mg1JgP7HfVEXAvNR2DAjd1G4puunFEwzfjdZHeDrEQPCPkKAVGS19/cZOUsM4s
31vkE89YC6uvthhn33hCV+85sdaf+IyyplQ2gjKKMzFSqLi65RTzjsQulT0FCpDVOoC5wNILLsRU
bvJQLuCx5qXn5oFm4K+wrPEt7FdiWwP76uh2d43mL6J5mEMsKyEyJaJOYAznhnc2ZSY6CoAIpJDP
ctGPglXs2NvFp2VRGHKB0LJmfNnufW/dbA4DBwNYK5lbJZhrsVE4fZYAhZwe2QoSVHM651p33mpa
lOvtVurD3RBTp4Wum3pGUhGf5H+vZyx76oHi/XJu64/PXti4rls7TPK94Opt4PEJ3iXVQmKHpE5u
UZ/SHxBuNrvY8vzGrCSMCL6ugcVuNgFAaDW213zDrEM9/lirUg51oPbkOyLp90zOWMNy57GXxX7a
CqRlxhcRMrpgHZSL/CbfpKcodE8NNuzKduXBu3ARCE/tgUVAJZA0xoVAd6LGjaPuo5SjW7aoYbtS
9B0B77pac5O+yowtd7GM8VM/mIizL0bcUvY0pRDFBY2mE41UbcoduupGiRHYUQKUEFqlo2fYqHGl
1eI26/BYi1VbCjMCZfEpaFpYCmR0L+cXnkIRW78HkSfkA2dVPWbGuXiLfYvB9nNYIgcSu5Mj9mAP
mxyODxS67yvDkhmvY0Hwry+NEv3M+srLNP1KYZhnNT01QgGHA6GWtER9wm5nqsz67zKXRm+rP8QB
GIH+Bz8czYUD3GjweVM7IRyiL01yjUk5sUiRj4XmAQm5GwHnXEp8MBEhdWEPW8cEolgk7/AT7KaO
bRBzYGGqUWAaO31tU7J0w8uIphu63/HQyN1/2+cyukg0n6NF3ykJHzSkIJZDfMBKfXiGkWkcsMoK
K6nXwW/TJv63AsC1c6FNNcTMcKy9fEnlFuCkza1p0z4LUJPF95Yqv1n8Pn5kcD/u13CPoQIsXFeQ
Y9wWPH9d9BR1np/82cTxjY3vIxr2pCFHOz0gLC8VTo7AAGgnVCp7RIpNBO1kHQzm9Urq6F9Saq5E
dy0hKJwQ/D6qmO+dBbuF8H4O0aH6MGwSbKePZBIWvzgUilY8cBz8hERUteqfYYrzN4xX9Ic0lWBb
7WEnBRPgviSEMrcHfzWFX55G1C6A33Fv5rZhENs6yMJojShMoOLU3KrcDacHuT49r7rhDJJbV9qv
L6BY43iYTeGfhdRmt7x7yhvH3hkHBUW7uTNYOGx3CE7VHhj9gdktII+mpvr4CFlK4RqT5acmzLQi
wzgMUGvehIGLUkgvNp/QoGTXQeg5+VN0Z4ElOqOdR/KjNTs0R2Ube0lmmdOrtR28fJ6aTAwG5ceH
dtVA2KF+SZvI+LCzmFqVJzyGfkER48khyBsYnx8oPg5IaLdchyFtvcGs3SjaYvm24sQ7Hhi8hV9x
Uj01oK8u2PyCN6UAaYFoTrRMq8Nx5XOo1eGKQYdsFdutSdp/9Gz67ZbNiy4nZxE9fyCjqZVp6FWS
QJUPO/30s3ofL/HItvZfLRj6biWIi8422U8MzNFnLgfJGA3m55I8EJtpjTUeUFtkutDwqq8Avds5
60kcUBaWAszkfzuqdTNILNYqrIsBGalTREkvKwO1exol7VF4PDvN2vLnNV5MgB0FpSofVN14kIr5
VVpl+hNg3Pdf4YxNWFPywANa0xz3dUzpHpjBSKoCEhXJSAJOH/lNXCjtf48EybExxDafYKTlZqVv
kkqJuuabvG3YVg0Q8HFYgjOgESDcZcZdikTzI1vYIICmCJzkK1zYLku6r2GGYavvbXY4Lc7IrYLf
S41o/q8wjAfc9Mpk9XlTLIA36p3cxs18vCS6/jh1bFqo0R9ZpyEw9bpS1mx36w582gmWeZbZiNx5
06T+uzX/05A0t6JLbHjvr8iyu/Fatf0Pn8LqT266OKBiC7rIN8lXwbIRhxMlBao9KDl+piJLFekF
0HzKDhnZYYCKlA0w2OUDdZodQMtKsO6eQeK41VeUzq81G6cYHf0Dwr9YB4FxbxLcB4nGLuqMHRAM
BahjbsqANNNdoH2rlt1w8ZHRptKZh8bAjjtlxznAxv0RdN2cgHavDgzN7PVLI6cmf3S5zWmkCvsc
Dsyqp7yiqdf9WnYoXu4chZlT/5P0DjHu8DxBb0uvlE59FJXgAIdeU3lW/2Cxoxg1dbZZT4d+8tXk
NHsproCVVIK720zX/cFt311soHg+dflvtn9TYj/uORuXsU5bN/CrKgpXIveLNalgY1EQHqO898NI
b5CsMlkYdTVFADuZm0xtpbX8ESpxLJz1mbZTXhN6X87XLjyThsmWo66s1gloLQziKUYRl+ZWs3+O
si3sZrZ49QbzXK+Zo1ayhGUpcLRr5RfAQowqgc0ZICVNsDJQOn2iiEqVRDb8QJUQeud1lEa3pcy9
3YdrqSmyhpIJoBhhRrMLQmdKFNzATAhCqjv61cXP20tsdA3nwGLHfv0jZQZ0CoMi5KaQatAD60Hc
w0Z5PFAS4lglQ/pcGYynZ58vHBMKXU+myeVnHptZ2bLAhhnQEgItSyEShlwusSfevXfa4a0CPq/h
enV5DvinWJii4A8mZeKmjYJI+xIeV7pkW+2alE/+qP1XAVP6D2uuAKPrYTUQp0iyzV4S6kFllRRO
yiwDCZNENa8Zg3FG9tI4111gIzbV0haPyaYmVtgMgTyfOembOf1wad2pJ54cCV1K/W3WokPeQtUE
HQEColgr9dERFiVsz9N4QHQK3DhcAvH0ercmP2NYBrpgv5EJvNCpLluhl5KZDX2N+70R75tHFay9
VNVA2T0z69X1H7M8lbfxSqqREU229t3WkynTeeBOpe27pVmVFRP6BKe5D5rDL6Shu88PspoPClxN
EWuu0cFHXPEfE2mSvWCrQwvnoYPvVPOT+dh1Eb5Sc/vXAaVWMHdbZHJ9MsaXXxEIlWbdzuy+6CeG
EDlT6ocg8j5ws1oTaQpT6MuFJBCzfzQWno3UmlCQguIdvAmz8ES+BdCNhlNgx2aLhuDuvxWy/LAu
8Xv12uoC+wMbFioPjXBeyHZv9GHWDFKNdaZ2ddKHv5bued3RhWBKI9UFcX2+OtAQh4gZm+WGBmaR
zWatDmCOzG1vnyrO8xBiDXEkMC5gLSQdWSOVIE0FZWv+0ONJK9qqi3qR90Rci+4ES6FSwuZYQkDs
v00w5ba3sHSY+8mQCZIu/9NcCWSjcpzyUX67SOGfaPIuQWwaqLIue+MgFIi6oz2c8SrCJ7j8LRcY
h+E460v8IfjHSx3MP0gCVcww+LVr1hl10R9cgA2Tk84mbI7lpI8CJDWkO6igf/J/tp4MIkfEWrlO
SQO4uqyKr1S/adnjU15GjtMS6WroX0ErQglcsUHkWlVGedeE30BUwgn7oGrv8WVdAD5ChQAuD4xW
f2ktrcMDs3NCp9xSGRv07zJc7na3hpGDMFaVylLFcUfh25vmUV9Co7yDnAP8yp6tQWnsABbuBMN9
irct/hZ6398KIEJwwD5CBJd1UyGVM8ifQR1tBmuVMRMHjlUFW0FfPzj76J+LPliJ0hNaNyr9sxJ9
PRQgz2D4ptUZF0VrVDlHkUYshHEqSswVjxWROUCPZ/hB/rCGVqWMI/rGHGYVIYdoGvEMHp4BzdnD
DSycazNeiRPRUUhhVXWHillcQBtND6O+JQ2/AUTZhWR9cgfzP3DTnqXCz2aKl847XgZ8nxJZJp87
+zIcybYx+Cw0g2JPe+knoBLiid9p2vpIjONwpnJ0r+9UGh36r72h9JWq+LPjU+hKEv8TLiBtC1ll
0FEoIOem5kakidDlX4MLL9omxqH31++M/M6KE/FtJ4q686RIR4F97Uu3cfjTvyqWTPCbhENT2g8l
vjHPOvtyZqn4x2+8zPQ/o4ohXTtEnq2RSkWlazle4ggsAFJXVcySlpNZHYIdZ88PKW08ZKl4pypC
/ZfiwONTz235R4cBtxNC2+y/gsH7Cwb2W72koiNWb+exJ9nJysKMDC6SfEn+UKhZrlqK+dF6vOGA
rwWY4I4KOiA0pd460xq90uYKyoySuzbHoHMNu5eFefYGIG0oDFkl2vPBxXXX8vLpUOdFL43gEQgI
68wIVPzWHlJTMMnWWuMlCR986jfR7PsvyInfDUCKtA1T+keuElKQe9oFsm2XnZEPF72y0oo4pKSb
LTaAAtQBg23gM1dVf2pMZgO5Jkvw2uo8mA2TdQ5VabfnqAO1JsCEI7ZmqT0tdzjEajU7rgarKrl5
MorYRWcISv/QIsGXPlQ3ADYtEqZN80JIjT0QQ6+HofihaSo7B8PguS2Hi1ZRb4GzsuLefxZJzQME
0zPZB+fFE3IMCuU5UuyIF7WykkRG0ERy55mE6tklKJr46VYASZZc+kHOTjJy3BbnsavPOuFgJp0D
oxyY+tOnltSEMRt98KIJMWcFIitQGFUaulbaXajLiUAv8g/Fh3CYso+jRzlgqUcP2c9KSi/6/jFP
/In3dqTaxzWPwBnyF+7KU4ALVZJBIyI4ScS/nH4smVzD0NFiL33FdYABUgdibkgr8Zxrk6bU09vA
QeBzp/kdnRwycP0OCEsELCkXau6sACMWkYWoj4njrV5P6KdYncCmoBd3sltN+AD4h13jhqbyYOnf
oCJXzMl/tPoWCrigFp85Mt61et/vO07TBk17jDoFKVTrNzLx3toTyKHx71EpPBa3d9SZsjt40NEb
851N75TDeINJvU3Us0jfC4EsvaS0ApiNvctNUIWXZ1beI2x2DwI2K8aeT8V9DiF5dnjcmsVlx3UX
KnSY4EqaY7cviiAjVjhq2U9PC2AcvMDU6BiHSOtryhoUc69EQ2EMmrSLIv6kqi+xk7UB3VZHohSY
rj4HYYhLyOVdeX6+rpC57oiTFXm+ipCfCR0icJ4sGGr250I+CfzU4rfMoIVEjOqRciwSgILY2dbG
Ws8zOEDlxvNUerykBV/Z2mBmaO4vwC8mi+jFeSPLj/t6MIWwXcBYblpq46Yv1xjNnlY2NmBb0YGO
q1xpmV3zArvm7EMs+GjDdQ6a3rEN0sW+Y9KjR13tV5UdqqdvDKXrL2rceYmQCHnpfJr5pSenvnhH
CEV8j3YT8zT3yvP2dImheFp6h9TugdEcEJAqgArFHVYg2GutLPmaq0uW4tegueZuQLVX0Xz6U+Qm
FD1oe7AC0ugL2Er3Qz/K/jBH3okj8aWvvqyASW3OP14INDxPCSM03dbme7Xw/ER/+7uHMlSmCsWp
sS+nLyyrFjFcD09w1IVY3Jn3smQpCKzo9XdBAI7QT6OkxekucpnHhF/KmToCe0wkKHxvUBYLd96b
PWKIC3HJXB9d7Ldt16NHv/SPROzsccjGtss0mJ1zWaONvyfA6eRspswJDheS0zrk5nYH0TtKuWCJ
fTcAO8rPRcSiC5FIbT5hRAxZGUTZWqCYUITtSmUXSlCCMwEsjODpLA92oYFKmX9R53JWRXpSvqT7
NZMVam0vPKAGsIxGa96vGFs5jM5py2zbUXMnCziecAtpMQV7wfBuE6hY32fXefakkv0AZ6KTgqT4
xlgQcmW+TDESPpHUzsWx4+6WJatiQTyM0VzNb+ay15h/+0PGrF3hG33pSeIAwreUZrvDNlqOUNin
YLuRHATH0ZAsiHdYSVPGQMySjW4x5FTE4yj/Yn9Zwuw4TVAFjeuxHHYjya1+2jAG13I4GONJzuqz
uiFcRObFYLcMfmiCwGOKKreUzOAU3yA7zgYx9Z+dwHvgEm7B34USe9WKW+FPf8qsv5AkubwfJFpw
10oBsJmtrpk0mWT1pt4z5d2B9nbk1mVpJqJQUHeDqj+3FeQ00gzbXlY3/NVI6BglNNWNG5Hhxa+0
3N3jl+1GhkWZvePah8HCPtPXo0OkOXV1nzIlFM200RiGOCUg4ppPYeQPuH/Porl5HMSPOOE3mfE0
ZbPJDxeSnrqOsBvhpZpix5U0bdTV5buo9xTpkMBF3QkDlY1lsVhecApDykB7n0lyPtBqegurzwz/
TU4pKaG3VbFkkn59X98UZWelZiPgPsVszmFX+uG+wD7A0Z077c+PzqQSDtII3UFnjFQfEMhapeQg
s/ZZ8uTOAQ4v6oiJGOUyZ5joUFLANQoyAt45H27HyDk17CPpY9WSQQw68o+Sftx9ulJ9H6fRNvI+
LPQY3Z6X1px1xVHx3Khnc3ezy9xm3Lfy7p4LCzgI9FCHtTPdLIbYVAIKiD7MSG4Pyvg53xXuKLej
xzANT7yP8yNp3S2T+XgZNXDUN7VFao28Ag6I7y17lAeToMDEYsoK9QPP5JPDKst5ymnhFzBkQ455
bA9ErEhdaLZZVRrKwFe9lmj2ywVXzOZXmU3BDXz1Dr0B19Mp4R6bIAK5WuA6IKbpquMz/tLUrjx/
fVWs2cUN/x+RbWMSjYxJ7/aBMm94j+CNRdkfZ8wkYVGHi7jKlgie0UdX1ESU3JWtVIo+Eh2PlCeE
DE7wGpoBdqfhipiIx3wedPJQrksmi0gqzCNkpgP7oorGkhbgsqMTVk42pfqA7P4CIGBwhpNUgs6x
p3wI5oGhtOiLu+bAZ3CBD09izsHds+9wb4LHDdcc+iakSTWbxhuSWaU7woTR4MPbuWXgpHCnkJ+/
5pNrNyrcV+H/a+5ZdRSwQYSbkcu8EEGQPesvizLfAfGE0RmpNAoWuSe8LQHioBP+xTgwf5xa6Jbx
MqM+XIm0vDly+bNQJnFAKsgAZ7S4/QlRofM5rgoKBIzPJEgTJ0VEsIc168X+yMJ+Mpi8umFSidYn
+UisWZTFa+nSPhleUVFcHqxevPMKHHFVr8scWIicm0xLiXSEePn8Xhx/0rENG7RYp4NTGCvf0o/Y
SuGt5xXeegeXsj0k9GSw/TxUs2rw286W5WTM5QF2gbL/+8soecwUNCMMW9Ww1pOoGZGLgBGKLcPw
pj6+ZuEWaykz1uvM417ZWABaWc60nZjgZSvQnbjkInf2cHWerP3tES8t9Ze3ITUjUqnBCaIFjEN+
bBVbECHOj0l0TOmFJaLHZKPvSClHKlU1qn24b5FLdXzRc81bRe/qp3QELCiOzjB5v3o9xVdvUNFP
aWBsfp1kLqYtPXbWXAQsuxbWqkoWuP5fn6f6YDmBoIRkalBMYmy9X3K4hodv95R3dJ7OFH22VkBn
WFESLb5G+/+VtcUVUzP1VNv9GLezTYOLXM4fAA8pFV1K5kjGDEIexxQiYnhzmGKQ+Vm5ZgLRe9up
hBXv7wbZY7besdhkA6ux4qzUugrAxDPX6mF66a+Cu1QPjcMZx550+o5PUqsFejirmax7qpYetZ0i
O5/qWfi7PEiPO+sOVxhoc208iUJ3eL9DMpBNcPHNIULmNx4NvnlBUrlN6ZINsLVuSJRrBemenVod
F37+mdsTE+s318aACWix7nEvSM7JzhBmqRyWOUGVxoutF/6gd6O9gXSgz7M+PzKagCvnQX4wqk53
lqOxYatRvmM1n1062IZGLqKguoMVUeO/gbQuyEBAy5Rgv8wztkEnEFZ70MhwKhkwjukMry3nW744
02ZvqHMepCv09jprmbPYPEFRXLdLBoXmOb9C8UH+LuAI3rRiBUJLfNyX0jEw5vjcymFz095WIUqO
rixSKKN7KAiL/xnnr+g36xtlHN91bgmnWAZKNOVF57/U3PnUPmgnWSax4t9JXVmDn2bWexUB0qH9
JL/4BuYdM8Qp0vEA4QrfYf2I10afDbqkb+vrYARXuIgKHpFDJQD7Qqp7KBFilnujXmsFXTo9ILX4
4gUUy1vOfq6NBBMQK6we251qLg6zmnU3hTKOzZuSMnHOxH13gb5sYCeo20INqI8Tcdt+dcusKk7q
MUdAdb5pr48j3/pdzSru/SU2Eh2BDkSSzB4bWCFOqtaw1pjP6s/cnqgbpAhJC/+M8Zd2+EzMdS6C
YiZwdgakVHBIQA92OhAe56I/ps7kKFLqYecp0MFmSvRPHaKVsZMTATETr1rCefRd2eDspekPn9sz
h30YslUleK20zOIi7HowM7aDFgON8m3vpoyYNblOr3Hz4JXVm5O0JMED+qb+kfxS7gQAKNPhJfPS
BWeV4+Sup1E5tQz0XkYfNLpuH8JH8k4o1sVNzKXm8kkCLIyPn7dGNG1Tl/3leRQK7sQcReYAjgCe
AZznhN+EHKgnXm2ZuBP3Xqs4LPqpgX1w5ZA0jPgcG4/noL+xB4rHg1dhib4xXHmrv/7AGMYY1fM0
ZmVms45N3Iv0/Fp+5F+cYsYa7WcSsJppqqKqk1eM3SrI8XEXM0zAqraYJUFVBkHeAN9cT6GurAlK
PwqCcgA89gIEZntyGKFjgFbb7YszX5S5RLv+pPOZq5ayZr9c5lglT3+rYFR8rXXRuf5ZS9pOe+rR
Bgw5+267mHIxsMV6wrIEIoPFtp76lCCL0/FiwAzZwn/E8KIn+xbTUPuhym0LV5bBNhtkeyB/hvfp
iXg66KsSAaoubUShcpb9F6U03CHySPgN7+g7XdDfppJPibLKnVbVhf3FjLMgeLTKJMh62Hm7KBtR
lXxlx4aw/zncGuNcyujvEKRp/+/ijWN4cEd+x9nBDuiuzJrUco1H1j08BdPCqwHXzPHVCHJMLd9X
prvJ8tr9dSvVD8aL9rxv0GdmVhcDl96XidPdOJfCLjdYhoKHL6SM1UBG1Sq9aHRN0wkyCqpSpUQ6
gYFJli0BCi+qowJkfdVjnnp+ICsJDmbRtgdfbt69tUIdZmkDMFJ+KZVWPAWm+to6xRnuUF9F9wXY
NXtahyWlIjifzHB9n8yMXqjMZgrkCQluvOVbeRkaOZDnf95vqe4q82sWF43T8ZeGKWjufN6mBgIU
TpzMSjU714EGeh+aPhk2eYXIKCdTjxkcWqgRqpfacBdMKzIrE5JPL9aSkyuK3lGffG33RQoKS8sJ
tiH8RB2h4x4xlPgTTYIDaS9lbKNEh5cNGMeYkubdQiDzA/4hmUmcUjrR5jCytkckHH8C7zd2NIVQ
dAb8si3qg7oOB0gcABYqUUbnb686ZkbNJeLd0fmDQB0XcX44l5pGpSHN2f3y/gVYZyxMlpYx1Mg/
Bm7MEnLTFYA1mMf8t04Wk0xi27v/+4OWxiyb4IIDLbfWTUDDQJkkW/v8pDA5EXLpXQ+9XMq9jGlX
WVi9MnVTIfMSzFbfujHxGuw0O2GHT0gvX/FCvJ8hraYJ7QLWzuHmCJoUj2nMgsi7eUW83Hodv5vR
cKIVqlcz1sww+uiZE6k+HvmBHaTvKSDX4Mpapndb3F54E6Jbj9dElLpG0oapk6TYhh4/ZO6b22IQ
OVWHSLje3dFR+XacloGfHS124XnSKyKogrJqaphyv3bf4SaTI9tus+U05rimvQ5FXCstd4at1H02
y/B8pQGWC3c83+oFvd2pT9hA/jftrqzmQpDOfHVyIWJxWP6EPx1WN0OxcgE4rENT7LTsh6eFE6MT
XPZyGbODdm5RXuDTigXYjanWtEVVfJ3H9bvaCBxkH5vba/F0uI/VFPc865F4uFSHEfojpJaXY23u
dwM8qZEMUo7/15WzObpchlQICQUvCn1IFI2qdWCTHtgVeUnxBg4OW7ATtepklGbX68/U6Wl4bKFO
PV50G1TopSrVDDwqAShIAu12rRKa2Lm23SufkCxZqkVvxmzn/0gNAUcriJptSpNgFKrByDj3yamX
s4GJYhUvDuMSzKyAmlHddQChMorBZnTqLKylGaS26lBGRorjDZKdN1b3HA/DqDVEEUcglacJJlAy
k4+GeuEacyfeAO3Wfl9OMOhGZJpe+FYHdWMbf2BzEovZaM9RvnKFx7+MY8kiDxxRC7077xGtVDtG
F3nVbIefM2FqmpeOkg6n2hd3rRHU/UEjOA9r0R+T4ijxDRmtyiDrJgW4p55Rw57oq4Nk+m0BIVRl
ci8zXQFKHIWykSDWg1cBIC7zjHpe+DNpbh597lx29f56Ydb+NiNnxHmq482HG71dHAgMKQNI2teJ
8oTa3nB8+TyX4IhHrHdoZEb9U4l0OhW1NxT/zpVCOIVEHuag8oju2z5HZgytkM20oYRE1kztv6/g
TuHysJC7+mmlDFYAUSQvE0ObtSLcEDbaYZz7q8lGDeGIClTM+tAyNiEWxHqGgPRhM0bMMDcq7eZQ
tFPJRUlsCB5V8fvc/AjbqHOWHFXhGHg1fO7rz/2BAWPkf/HczJMeC7nfZnGdvw82GhIhZpOQGfue
irXtsf4HpO/upC7Tw87gKqXvOWQ2snsEKgAND/O2SO8zqgPQd+uSP5wLR+rz+GbxuS1yuIypXeel
/Sia3qTMseV8BF22CzloE/FG0w4+nuCgSUdbWEvsO/Ywqgi88zt9RnlodZuxjA679HTgOoxlo5+Q
q6wokCZw4T/EFSLbh0qF41oGY7HekeKZaJYcVsVQrktLOF8PC3MicYJ1IJmC/fLxBSg9StdmjsU+
2aIL9Um+F1UXk6dWvyvsHjnwHhQ6s4q0HBn/GwBCcCE464tnS48/G0s37HflvVBKuviJsrnVWmrU
h+Vl8LKZ/8gmkg/gJDohEa0bZQpMbdd3SrvNdwTDSK/0jHJ8ag9WfB0/G07WmEHD5zSD9I/t/Ozk
r0hfZ6iOCoXM7JUZ8s6ekgyxrScMU4CzGBXBn3u/LNHNhv8SPHlU5cTcl6dCl+tI7LZbHh/+q5KT
YOGdkcDLkUqhdu2YPNwwYkDxMhoJtK6EKF5z/n0jUoYay2bp7FsoSH2Au/HbrAvwasT4obJmCsr6
5q5jLKyRbdMB56KenMT+LxyagS8z2Z8hoD2rECNWhIAZlR7sq0ung6lIsfQw56KjhlSV0aPs8BBf
p+HBufwjyH/46isO7/+ma7nRq5yZAK1TDf2v1Y0DXxUOqvDtAfRITIAV0Br0ptommIqgdwEH6gtr
IiOExnVZ0e65iVZf0yKRMbL0Q/NOKEjhfOVmvxvj4wnApq+Hq7CerziUv7kFtCVQbJu2oinXTFBk
iNCNUHHV7nw6gx2I6VdLbjCfHQF8XWQ3p4Kjc4VxDAsgEUFtfHLnhtHtSry2qVQnBSh6oeP5N6eu
36yL71vvTfPpC5timlsMdVfvYLAFLHQ7/wHGw0e6V+QGMGsg+RsL1IPuJ4quukuzkvTSXBqEeNDC
uzpdbEnVueaONQt5ew6FNTUr2cpmNy05W7nPb2YJMxoV1kL/0PSVfPzttWrL+Fw+noYAwoYpESMG
he1ZhALYPaFU56n5nKpmFitDsc5ilBW/gkD39Uar1HITf30+PB9bmYADAbfJ6PutVcp5a9LhwbL1
qpyDrrsblO13b84tLYmK/XtpIuMu/dXMpC9awmEWFhrTcVvspbMw4svSj1ZzKWeQuZTTR6DGnUKE
5fXKurZ2cc+oIOhP/0MTjzQJNDDyXVTQGK8hgr1deWyQaQHeyWFg1y32oBD5ibR1e9mTl7Wjgq4y
4coFVmGmgP751VgGAk1hiBIMQMFXdHKqJVjuDGL00jnHMveWELPqa2AHE68G3IoO7mH8ExbHFiXM
+f7lgjZGDyv3OFsj0jiSGLOLnRopguzbWnXX2hL2o+XDFOmtgtgjK9IH+uYJZiuCmS3CZ0Z99ppn
vpaHRl513wPGeOzG6O2cTOUTKHouzIMP/fuKRMvDTbxTesWW1ZB0Vr/Oaeu/ZUXhgzrgk8hUsKNO
t+bCJ21aYOLcX1JEzP2uWr2qaOIoa8FDol4o58rRteSrbK76J2Bp5EwbuMkbwZg/GOO5VayE6VCc
7dAjNwLvXaBOVWYeEgcZ47maF+PwwF+v2pDuXE3yeVl2WO7nSxql4Hj/L4Of0X5J8oazIlFNili8
gS+R4pyb5V5Avz7SD7cY7UCMSfivZTFriZmRlULj92cFw8A6LLiTOkar/j+UmsanGUXPaotNR5/B
gJf59kh0z7s5hWbHQcypz+oIjtG9JhZib57FzzaFCsqqymmN7JK058qF0L+OLux0IEpPaaeOFJaw
T7/HNyqNGL5pMK2yw4Zg7+dubrKTokZ+w2v/A0G715BsJ3aIYg6E6bxU6nKj6CM7vQTta3XU+7YE
j9m9bFM2bz51x61ZA/rp9q2kHauK3VOdxAWcqVeuL1tNb9xfPAKKWsiVgc9B6PZDGTiXdQV/pOZK
gatTPt32NYRXKu/y0fEiGyaUGB+buC4czJR3ABuB3pQQPT18S1T7HjKI/bgOqYum7s4S1wawOVqi
SYlsn6Xt/3xhNWMTUEK94Go8rrlaDbgK4/tiPe6J4yCVfGZZf2aqM7N7J9XUP5TseOyifE33FAk0
Awyt8ATiXIq1HPXTXb8fXYAjWaeREquTfbh2QimLn7CSFJr8CSzhwcSkFACdgUWYRP426fy1T5dN
H9vgdKyQbB0ATSn//UJgvsYWPpv7dmX7yIXLyP36DJalQuyiGAVlfIz9t0MB1vqwMM6dmR2V8FD2
/E+x+7HQ8835E+f3Y6dy8ADL0vBT9mB/V04HZdJRaGWmUWJVyFki6wvOjjiwkHtGn5wz8voep7Qn
vA2ebqJTo9hR4eWYZYshN8XklKoA/G4x/bjC5/bSWzh5Ic5/q11JbZXrYjQvmwry5O9ZfG4EcTQu
BPoQWnKSXsNe3918gmXOfkCIkmsmlqDH/vExyGrh4TcdvjDj8sk//1HgjX45bF8wDB16/kNwJE+K
yiipRP5LLMn+bOtCosB+ERv8v3El1r15yl0etQPZovqAQ0ph7CV3SqWIJdkSKUdR9FDyy/rS7kms
HwWgN/IiJQkQXEsreAbA5csHDNMZgygjUgow81eMJc07sKrTG/56qOkKQh/c62evBOiO8KhiBLbR
7a80DawxGFOvfeInml9xbaJ1xH3Zj6l8BfbzHiLz1wjjlWQC9BKyE3PAlpJMa6lxX8jMpfQxMIT5
M0Xp5zmAMWULbQuOiTMy1Qjwjtr1BG+66klfWpAZ809PUZAKZp0XSyZ8OvhTYvI1aQRZpyvjRq7E
ckQODfG0cu8clf0DAyCOpAOYuvtwUlJmwP9A8Nd701v1i1hSQtD8AasCkS6FXFqW05I37m+T3bem
hyIZeiY2zQQ4JQq3uta010iped1herRnwHKElNBQYu5kDVgHfkTBulQLlSXZUWYhon1EoSquXSgI
wfgsS0QNLiAZAuL9gPjWL03Eg8BVrXsnOD7PJ3zEO064KDZTbMB+yGBTq4Ekdbfytb2mfSTtaypP
Co+yzvERgTh7/tWtQPWzs1y9swYtyGKjbO2DzlSezRPYDN7yO0k4YGY0HQP8HiTy0ZRDbuRBoQBP
2ymfVbqPpkPyAY1UikfpzNnbvRLTfF/wxIp3uxn1a2cuEwoRwrRLdrHFB9KyDXoAhLJtSZno8BH9
/tVlwwiF+K5chiBrS0DzDHGq2c5L2QrYiULYz2K0hB9OuJ2xQGqv7oTmf2T8G2UP2X4sDBa39i1Z
EN9+cx+o3SzfEg2oFuix+21hTflvDGcAccG/LhYjzhXYwTe3Siwc5l68GVgycoJANXQiqOI1V33P
EvZSaefqgY0XrZLIVErH3ElJTT27LP9YkmUln7hQHFeNnadRnwlWFl6GUPZCBltOKd0kYlPLPiAd
5C2uaNoHjMM5TzkUrrpRzez1NAdUyu2KTcfEH7ZllSrM/TRoobj4GPBH/SyyChI/Ezu/4NDwPG8/
PkoAQFDZXKNDnNH/WdzdgnbO3b0+B42l21vfumveRssgEbBMZNsiBL663RKxO991tnK0m7ckxxm6
/aOnVVzfDPIXlyLna4I1FJue5SiAiUxwLoCPEolm6rbxMZxZdN+zeZQfN/xtEySeXWs9sO4F0ul1
effzivIA71GrwyslKTjidvRn45ZW2OduF1yxLcnwj7uBGOhfJYnv7933zhg/0YqGcGGGp6z0Rlun
GFpdXlYWXPIjZ9kgD6CuxA43esCX0jUP+DANKSQdBBtVepn99qiYR7fq+R1JTVV/Nm45qfj0Urlo
Z6KM3X2F5aEQVGpdA+cLlsXx78L4GEtkYr/yqqAmaO8u/bos058AYo4bKmOLXb0nVnxrbqK7xNj2
Tb3gFELzlrJaFYQjY/OQ7aL46heTnavzxm/2IxTw1/uNPX2D0xIjNKONL+adRmT5rCHRxqquqr7e
CGFD5OsF2guUG0tKpnBmCVJ4duV2YP8FDGba5b1KNPuiLinHecfwIuzo0S4yIT1yebb9lthJwwvC
fu8gHOWkkod30zZJBptj/bMI9pAOYXttclkTL2xeOEHIuXK+oZYHyPMp6uGuTKJ29Xn1/iEHtyne
yYsOZP7HB46n4o9TqQxK6h0eyM5yizoRfJRTi1XfvuSU66LINKchNT9qBSTX8GIWk9whDME94YWr
AqwGR9CeoXntxiVs3EIZyy+2SiZgkvSQZxi+hjazJ6ioB0aL5lPb61dqrhjeiv/IUx4pbIcmMkZ1
SMlfagqF28PVTaWjML6WBA2Y9Yk++MV/MwymUFN6LueaaqctCVpg9dohxo5DoMVP+EUkcFZDut6Y
4YIfhQx1kRiohTZJRbLOvO3rm9iaqjsBpSpBNiVVQES92/hKPeRyDDh4wlEmJo9UBJ+Cj4Sz6VaO
EmAuOi4nycB9ixuPolvqYMTGBM5ZVLEr2sENzxQRgT8+tZrpLjyIuH+YWm+S/+gtuwxepq9vh6g4
driYBQaJKkg1OKNyTmB7DXHawWcuhQRQsq8uU1IoiuaNzHv8RtXO9vBkM3+tURPt9YL1LLENe9y3
g6rBIjJ47DhHC8jL7vlP7WheuQKW6mfDCoIsxPkwvhb3iaz5B7stl6Vmz5mxKo0AfI0uhHeZI/40
0T6jLHYCeNojL+/c2iEQY3yXR6rl7YGHucjfVgQL5W3hfo/Sz3xPSgpRwUrz608Ignu3EBKFh+Rj
LEaFGwaQMLkwzg8sC20I2vJW9KAsFkZcaSIazg2Dna3IaSTgc3kLmuNH7tgKEnjnHo/Ko0KNLdAH
gtx25k5iWnicFRdBIPUUeeuhdK/9F0PytsLnoR7MJV4Rk9NVS6KEwp3G6dfBz1cV6QxAuG76u4/8
bnuW0vdRHfg7en9d6wxZQybpmC5JElq4S6ybRbdTG1G+hXxGAVBCXqwlhDh/4o5dYfe9AqMEr66/
UFYTl/EkYpwuLdkn7ydMlKdz4QrS8PIlTqxkYs2uU4twv7xcB1qrQEcdVXLMlr+ZwcffksngqYyu
RBGwI/d2uJ2J1HNTFT73vFVvjE4OjxC+fwgHFUflQ7rug0LYrfcU1/cMdEKkmLznhjQS5LcFm2US
P/pKLYw163lVeSGAHO6v1XAxMPywbA0/e3ktK87M2rWo3XHTyl0LRU9VGaJAh4sZnWfHi9RSEqxD
OQxaCz6nBXXGAiPxBbDCNDIPIvppAd5QrK0i3KtHulSGn/sTg4YZRH6RuQW7izZO5HFhMUjXX0Ua
GvjPVeBBcu+Aj48QkOjkjJO9zaMIxzNfBmEJIhAsNxnDxyT7WYFSGEbtohr/472/+i6TLhGL+T0b
lRjhWVtlGhg7D1zdj5Mamzvngp1LnRefJDphUR6jSQvVOGzolvqR8iogtBZiosgDPxNYsTuD005H
5hx6yDX5D0qv2AUiPmkx22aQxuPDJa2yUFF5dv6JZaMRrtC8/qlXQTHEeHqJqqaiEme47Yisa/T4
a+61MQXvJAhWWM0+jkYgvzjY3SVqEKdQPz2/4hV/IbfmbtAYEbCRFfeUlifDE5bxCcTQ8GEB0yub
lPiTWNvdnIB6uB9HloIdYeZfX2bVEPvmb7alCpzIOz35CGJsXhqNiJSeK9r+GNO6040lohz+9UTO
GK61JU1hVYNDovG10Pd6F7nR/tFICsuMK18dBX2E3KOn6n6/GF2wSgpeEIGEkT7eKhjOoZe7fpq1
K62qnQswtM90s+bdaAKiQcXXwkOGYdw1QfgU9qfYNMGDqGtiQqmX4QRLCOVgUloNzxCUnTaf7BCm
J9zrQAnszafVV1G73rprXSruJtdrVSsfnhOuYjtIC78doEtStCAnZkFxAv6vgVFOkofzvqJpyJiA
fjq3gjkzwi7ixqEVfJVVUECYEGp3vGoSFcQtRKSrTYuvTNuBs8AUhLZLSLTMp2HamfwUFvs/k3WC
VF0DaZrv+ZdEfCimIwt4JtecDG38N6OVhCMxvCLkbeKlPZJQqQNXzhkxvo72dabEy2Rr9wKpYb68
bO60UCsDJVPreJxSl+eOpG9CBAeDRezXCXp9ch5BvVPSPmYOVh1Plf10FsxOcOoPuW09/AYwJdUu
q2vOLWkLJKwde9AzShyQvCMQ4+kwC1qq3bowazI5v3dpTNWDrsyE3ZUXpJc8xggU3xjTqApXcecR
cEQJ3xFs614e/6bpwwhM7gfSBCiDxtp39RqYbVU8cAvbHUdCRFrRf59oKPfz19MEyNB/+hp06DRm
p4XWaU3xV9EKS0E4+DLbbUyTLgihOBxvl5797fpnNNtbAD9w1lCStM/VIfOpC3fPwjPObL0aixa5
0X7TO3fbPmqRFSDzoHJpxhcpD8Z+77O/vPr5HS69MC6tgVv8uwuhEcW7DnzaSv5Rn/0/vu8XBj0L
JmtviMSq1PMT6sm/xsLQimWLYQp1p8/LLjA/fwkMwYxtyY90/JYbBYAoPzKuOlfH+kFwYy7IsXuX
70PUCNg3rhRpF2hQACtkOjjbV6NoGxNQDZZYd0wVZ6lx8A7T34bw+ae8g5+OUJ8BsN1+oYDwtLTp
8kmkzoWXG5mLmVZrtWIxVFlF8bRO3Sr5Ow4WbnPFLAjlxcYHfxlpMzJdC//Q49sUGL7xzrg5Zg6h
Pcr0vl3V2+gr29tn0a4WfnewbeSYBWuHVhJwz5hxDTMoXCeUXmEMSlhtPrA1MFYxGsMFn4aTH2yR
O6hirkLLlXTBOjf7+nhQ3NYXbYrVg5XhKcb0CmdGmxkvmeaCT37KngAzy6enTmQiPfaIsAaBmnPK
+5sNYsg0O1asGqzkP+RNkcMO9OcC+niVJy5kvDR4mLap+HJWE2LjwBcxjEEPGa/5vytrao5hC4Ul
cqelr2Pf/9+2KxXU+2Uc7hbbAzy0kXddQNY9sdaA5bkZ2CWl1TEKatdCuD5vzELVqdBXmguJHxXP
0kGwyWy7kg9TfEz1Y7eQ1b+9uf108TB+QbGRPP5tV6xnccXci/YrqQZs9qpMdTVJgG83hCXEU55p
ueNzPvCOhxG3lbKFTmfiya3P5H0n+oEJFImdE2GT8HGkzfjPPwTcJ/yFI/xz/+THChV1LrGjl709
eZF0BX2NKosx+SzZDUZdaY88m1p0c5kurRcweT5YOHc1h2yEV5K53q6IEjteUXTH3LBSJ0YfHcQ7
njpcldtR8s5DlP5ulZ/2iJrZAheXFKDsKr3Xs7uo30GqB1mZZ2dFNgJnJYAhznRYWCaPt0dwCdRZ
PBP4qq8ajI01u4nW29s2MoTINR/g01I1CHQ0eygc9hj8Q/fzTA3l8031r74RpBNkktAt1KTyD35t
ELxzGJV6lphJsED8pZnTHFwYDi9Z4N5MQEr8APlF5oe0KTVC1rvJKC1/NOfbNOIX90qH5gmReNmc
nZNEo2ccwTqALm/0id62czeOFW7ZY2X7ppZwU4qBtlA0rgJgmMaKvX9tP8F3wobUFJCt7xqgDFoi
KcohWttNeefRWByo4jxf9hk1KZAVCxDpmD2cICGb5q1OTakNgCrjcyUPZTtFQTgRxW++UPjMk+St
BVQZ5uk2cj5g9KIY8txdKy1t+xnsDDHXLnaVm8wMwLOAHuQcmpL83MsvxUaqFPOIhRXjIYFUakW7
6iZcZJrgiJpZq1rxXTrDhRyHz3r7YWq9iocvXTcg8ny6NASUEpRGDyGE7Fp5RjK++aZ51fTWmD84
zSEF8eBf99RYN8XNxPg5YWvn5LUBBtLQpygqOSd4YdLAKwSrp5MGeOfJJd9S3svokkBroJMu50fp
Si9lxXbwozkbVDy2dyprhAZ3wSV9bipttaZBpIYjUKw6u0/QBgVki5lEytXzjyC/WHDL8hg2QKM4
xk1xrhFjflu3B78adXHPWTthyTZNm0RpH7HfMgSAr4FatKtsZgweGtCI0wHDP46uMwmJjVTcecqh
XGRhhoCvyLB2jYcqi9gWQVIvVzNS+0C2vuN+1LZ9EbZL4CpsSeG7w1RD8eCbOq6buMdGUNjT4kW2
97nSo8OpMdvr0yNPYeB7/NGMVSR+2AwGiYiRdqodsYE9T/IRgxywqCo8HhYhTakuVApI5Lz6aIXn
pq76ObDTyMKQKs3npNCJKfqQRwEBPTL7bp4S1zxFPqHE2NkgmZwWjMzsGbZ7iEfhjFvUVIP5hImd
qmhBW6Soth7cXVPSkvj5p7dwTz88sIlIPZGCwR2AhR+KN+PjGROXEtqlKRaPX6Z06lQWxmRUbrKK
+WnETCw1doxmPLCuGDSUwK/3mmlzuLlVXRdtHenX7ri7JNpsoz5IW0ml1Ofns6uihUkop3EqUpiP
rXlacxYyanWR83fxaZ6RtLt5ta6xAf6OjEDS9H6kZ76Jmzm8+TEf5Vl7fxj+bjdmwTHWMRxH3p+j
M3WpEyYQQ5tjei0JBjDqoRihCtANuDclH0s/kyQdAGgOleEM4hsWFAX5zWd4x2EAsdxCCsyvwWlq
GnXGfGWSsXiR1KWYe/nmvpykINUB/jFnoS8h/TYA8Yd6HyJfg1gLQos4ihFXbSRipDeEYiKElNES
fZnbyScMSazCsdqtfXB2WS/8jBRbiqXEPdUVN/6Q0dxzecjGQF3BB2pDpHaNjGQQR6mWlC9KgJI4
rYFt08M7EoZIJjSUo9nQ/oQio+FBRkrmnrz+G47vX/2C19AvG8FjMga0YI2hnAl0X8idTtrtSMV5
DGlte/DOMuAKgR3sM2QG5BbjD5xV2pNRvO7p74wKndkQwCDHHOgL+hhK6QVqBKRL5Xk9DHa8XAMI
ixP5N2Ny3wS/MFycm0SFpD5JNnXnVS90OyzfIbpBTUziFLYEOIVG/trtvxA6N2XIxQPX4zI5lhqI
3WyB3ifgUbisiM/nPPy9EZgzh/4SaACZVYkLxfvGbezFbwfvRnCMnnKFAbCju05bULVI9cTxTI8f
afyuzEIrL1Er7QGn1RtMSUvo/EtXUfhLqsLguxFNRso4eVr9IJ9YrYIZbLln8wUqYVARsFFNLCTq
K/wNWbFexXn6sgomGc5esfNNDigSOspLdVhzIFhqdtks9fz55gKHXK3gbw0OT/cx280e/h6gtSr/
3klVihvUw7ueftFwQFR/Semhop19e5ESL6wjhkRW/eddNESn50XJAGmHHVhER0PFu6+5ZcC5u+Ry
thRDQYdST1Bk2vB7WqOfRnPgmScR3kVd3V5Wo0tbFW4uXMF8ugm6OocXEe+Sk0tpqOqM1F0N3Vxt
LhHvhB+KWHG1NIrShBdczWGYT6Qy4VxDydSLO6XLVfcdSjLZv1dcTRbsj0XNjyGJVFKo1DBJkGsU
UNXGHPNF3PS0r00oymYf2X+FsnmL+Xpu2+7bXloLYXJtk4tLTr5Oltshn4LucTKIo8IMjCQldaNe
+GjzmmB8/zBMouKYN4fVWB5mi7qwJ2mbCgqeILGnL1P1UiSV/pgprRFMHrMXSAlX3FXG6ZtmY7Sq
P9mVbsAPrHbuvT2owpTRdmdfyqczcrlXSeEVYJJa6+KxzIjemjFhrv70zNsgDd7prLeFHJeAmoRP
LdRqpjMZz/EruCibpkCMizCiqOUkwFWcqybzaQe/gOFZa12850AHRo1f0q4aqFkex3YAbyxG8xnY
HQiboBUTusetumLwkEhOOPipbrN4sqqjcHFDdr87TUbNdMKjxiwYgW4Lfg76S42RbyOH6xVUSWAt
YkK8/Fx3zR33XCJ9qRti2ahC0V70UbSQCiqalO/SzOypjN6yK2PJzDvGbIjrhX3lEYDkYpgPUvPc
9a8XB6boalPJRpXXApjoDh0MrzLYWv22buDqj7xf4AsWBKHpPaioMVoof6ELyB9BAN7Yxxkqdjxk
azMQskLxHfVvivEBuV3WB9hnD243VO7lkKnrbU9oIl1f4oVzIijOTJ9dCsP2F9ZOVj88GLto3e1J
XnDHu2i8UuIXujTk/8yolrS901jCUS8KAml7zv5AngIwXqgBH/jgu4oqJgUZ1Cf96j60MJZbLyPp
CEXUYfs7KcFfhiPG0Mg+0r7Z5tID2YLFVF+oleleduGj/N1dcEY6kXtFX+OD0IQ8eL0G2m2vWa3z
bu9eC/BvLPxgXjYXIKXDBceM4p+bYxHpN4/ABOpRk5NbOUoCujF+1/kQAO9f6m4UWWZsRcKAymrM
R2ndd/meXDK8YAxfQEBnoMWPjU9qKpjhfHG0HUKgnRIGyLfZmDEZigW70t7HuL6kRBCZ1XjNSL9G
hTgkNXbWQOpjH2N7++nA0i9UaUMwyyPJECp+r8hY/hCmhHoGo9hz9s/wnOHhlFUpZMchqUGd8vxa
4XnArPsp4KQgkVs9TBDQjdhnBoqICU7ZfoOWXguNnE+r7RqIzlF3NR+B9xuL411OSMqAOq3wXpjZ
tdtv1kEqyMZmp5NRBP1my2DyCgboxBAVVkOTBMIMo0OUdoxtNrVGNErn5Hegw5QaWd1UdfipnKeY
aN2dtT1bavJxoAu2u2rSaiSp202BjLj4WmieMloyAAhs36heuqAc8p1SDj9+f1XkfdzB/aR4KAHl
/lXbHJoMiMsZXDIwqA+HG1GCnLZtd/1zy8HBdu/S0azgJAgc/2i+sZBx3yApBiHwem3NbInW68te
3nQVNxW1IsMWojqyfxYQcqXiL/Bmoe+/vtOCPTlJEnwNLjjnzkxDN+uVFL1mc9iJtyJ7K2L9UAqy
6oyKJDhqbN0freCxu/S0gFTYSsUHTq3f4e0F4HnZZniwbarMVP10MueHE9s08dZRHMNfC0qJBA6m
NBwmuLVuyRA4GcSHHKH/zfTK9lh0EB3XMoeDc6foQw/0e54OAM/hZU+dCCgHJM3cFnEIYyzsNlED
9HDMDpV9mZ9cb/O1WZWgHO8txdPfFskYKLivmAKbjDeDhSQT6hFAfsDqP86tFD8s2lEYRoZtBDsX
SF5FQffxJS7BkXI69m617XwyNDjsJp8lrTw94sxTqryijzWeJC7viCA3T0+BkOGkofs8OrRvMO+T
zFM/DxNR7RO+i51HKYTPYWWdDPaJUpsjK3KpI5XEkFklpPPqpzxAv2kjZusSu9fABdzkqezP5+g0
60nUPUGPSAQkD3uW+uMWewDpLRbbo2XixFvX108L7ySBO9C3nwZuT70LIbJn8CxAo1PT9ckpjKCb
PwQsYGwKaWeUZQVwTK26ItfJ4Qg3DpIGjpY53vlCaA9byyAaG6izA4JsoPuF8Ij9zfyf6eMQblQI
NkSTgDLOxue0Qe3bz0Jm181/vkv7PpLvaRPk0ht3IlS8Ycy1iOoiHfNw9wxyWKo+2FHK0hdwmifZ
K93iqMkrS55oBEA7rKYzidE8O2ExTery2AEWezPfh4H9AL7mv8bVmBK1VSlTA9mFLf6vEgh098uh
zA46IwEJ7ujYuI+UxvM3T+9pVvpeuXAEYXFFCTYJ+wFQ9zCa2WL8buxk7JQh1/bDcsZjTLRJU3Hy
x+PWXMFGVl3Ep/fouJMMCtynecPHL9qkUtsWoghbTFz2+z7sB5VaPEusITFOoleZn/Ktnn4kXvle
lSq8axZfIEph/kxLij4A293SFhUJR38q0G4APbwzx4up6lAOrBjZwpllSROKiaD4p9v3RUYqHbuA
vlJAtf6SFRWU03YKuT1CA6kCdgZwvEUGGcC+u2CCT8Vo2+c+Wd53EMiNWMGxG1HjHp0r9PP+qNa2
qFqCPAYwrTO2+1g352d4avJMZEyY5k5ty4LrsxBo1V3sd88UHk2VOZPGjYiIL+zUmrAtQx1sl2jG
YiVLfPNwv/MQ/TktOo97LclVSFGAVYd0OhHoB0UNh+J5KxhFZ1hnvPKp4jHOUyxzTFpK4zsVy5wc
NaRFlCzO7IvFf/C2GT+joslHKZlAdlVDdh15aFRBSaEPT6TucItkC8od4PnB6v1sEbznylVPgzvp
qOz6cSl+P2E0uvLACxjFdKNya1y5m77w4ptFPn4QcZXmwEXVAr2AkmNPmKkyzwVY/WvK9gfhR3Tb
+BQXTgYrYaVyNQ2B59I+UF2ElGiLgziGH/yMHshSPUbxbsGXnIHyQVXq5MLyINUy6Q6uWfxJHLfX
vaaqEQZB6jhLAskY1i/MEFf14QuvhuzrP4n5CBCxBzuGDEZLBDq5iFt70WeZCTD93xLQJ5Dq1siC
UNEH++WdFwqErzHkDgsUjWdn57I8dBN7d1fWVA0mah1sbxwcAf873iZhbCUsmI4HLWQnHxpYZuP8
7WAHLNa7vi/75JPvr9c5PcZ5diqY1+k0AaN9zl9npra4lSBbrE7YxY9Lqu/aH+8XYExsO/RgCxQx
ZgrIVz857KnhfT6ulHkcOIfvcTn5FhLN6bF7ip/8mXybAvdsnRRpCzwfQQuKY0r6UcdyTSXlX4LR
lVw7NkxakmhAs0JCo1+/IO/6G2L+ThKSdh/9CxuNUDfFwqG8SZFec+1MBxpdeLAy/xid8teUOnAH
4YmcAGvrL67Ql1OBo9NvrFWqRQRPQEZaQRTHiQVYQGdoHJ9ROb1/3Ct7yV6Xes8Ss21CZe3tIje3
xZ/TzGlv82U2Otr0vYev8wv8IfVv/wH/PS5eorG6o3jsjkFivNqJ13lk/FYvS0P1EfsHMyD8BplX
ijhsuMg2UrHzqHk+Qaj96d02xYymkhM73Hn3lQ8EU9kh3fEz3umv8DzVoZ3GHw9Gpv5g5ipp8VCr
xGxUA3tjjjD/w0vwV6w2I+FUmXmrIi9cPRpVT0Kmn0rFCrG1ePC31hTJ4mnKVjHs53yKKbFxEYHT
TuDrTXDqLt0XhCsOnwgsEMw0Mem0EZz2FldBtEk9sp4UwU9ACHqKuCJBNWtQdgofGNJU+7tdgN82
EnajDAj7GKO/yFgxY1WdzSy6L5XF7CZNlL0RoAWPLLlJh3fU4c1GlkfsfER22EOLihgSaAdgakbI
R1zp4JqYIEzlhYShKz4Md0Dk3mLd4bRfGES5iWK/peR+QyA3mGREbDDixIoFf9+lUF/ZeQiXzRoM
AZ37NemgakO+8CkgtPY3Fn7c/muvtPUNifdwziuEdGDXEm8M+uYPJIxDHOnbC5KTKdGBYSpDV47e
wWWYtIj3+GgzUxI/6fnx6X3IyllS2e+Nrv7YFon1VmkQoquvSdzLza3Pu2KPULd1KvAF+xmCVTRg
JWGRo2bf76ektK3mlYH3IKprnpJ0WHGu6iGPCCK0Ig1/DouX8L/ai2SArbVb87q3+Qn5CRQmkysY
3Db+Lntd2oZo0pEWI3Kbn8699HGQaDATde7ZUCJ5KvTWzSQ+pDqQMvYkf39HPhUlcF55LOZu4eHs
tXkz8vQcdc6r/GrTt4XdeTtf0FBdW5mGMRuDqVm5AHBxYxWZBCfmrF91GA4xbpOVd+PlckmFpNMI
LmUqlro1vyrCfsEoM1mnmgnNRY7tqmJOwqlHhJe16AY0y/XDJhjCVB94/yFnxAJTIkVH5BReetoM
vhPMqLGOmY2qKN2fvfjkCSrOtfl4b51960LbAEXyKwmeObmw9CmRDgPfeZPclwxDzh13ChgPRO3W
u7eeNNIKDvmxaXrlJBVtwhDhNQy1uQm7VEA+/EQ/Tfj3uOhMGm2fM2+56R7zeG41F+DfodLFOlS1
ciySdmM28x2rtwRyU8szqk0yRqUdt9Ak8tqR3XM5mfRosEfTXBw8ocYVq/XYOEZgKUT4NcdGvMRS
f44kqlmqYCCVKXZgOp44ywE2NdW4DvWx5WaX5aY1thkQrMJKvTKGgGrtPE8a+jwIpiCC6pvxRAy5
ooCCHu+XahBsAKz6m/r0+RAdsHX9Op3CZICfHHbqqoHA7RAxUEbMGaV37cI1V0MQ2O1Bn/ezjkJc
CMYl13sPT28PrBl3pN8AwWbOKgC4LDuTqQrqLw9etcYJ3h16VEy68o0ucT95O3cJda7qO6whNgu1
9p/fVCBOGkmuNS2nlKuBcDWkOWUidUf8iNRS+Vfbzyed8El9IC/blqIpEK8eTrVp5teHxs+FUh+m
OSXbDmjoz1eFrynmEiFr+6uqA2RduCQbcMyYxP6fueXLTnug1lMdV7hdgNujwkJVI+Z2I6OlZFhP
N2MplLg7WK0mpRwtDGEDKZXMXnO+tk385syaUNWpl3F94xaBUWFeHPI0napfoFSOa06Pcu/RQ+XK
YdUQg9uBgoCZTc6CUI4MgU3t8CMV1F4tjbsT7hgF12T/b1c+y+YGa9Y=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library synplify;
use synplify.components.all;
library gw1ns;
use gw1ns.components.all;

entity Gowin_EMPU_Top is
port(
  sys_clk :  in std_logic;
  gpio :  inout std_logic_vector(15 downto 0);
  scl :  inout std_logic;
  sda :  inout std_logic;
  reset_n :  in std_logic);
end Gowin_EMPU_Top;
architecture beh of Gowin_EMPU_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~Gowin_EMPU.Gowin_EMPU_Top\
port(
  reset_n: in std_logic;
  sys_clk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  scl: inout std_logic;
  sda: inout std_logic;
  gpio : inout std_logic_vector(15 downto 0));
end component;
begin
GND_s9: GND
port map (
  G => GND_0);
VCC_s10: VCC
port map (
  V => VCC_0);
Gowin_EMPU_inst: \~Gowin_EMPU.Gowin_EMPU_Top\
port map(
  reset_n => reset_n,
  sys_clk => sys_clk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  scl => scl,
  sda => sda,
  gpio(15 downto 0) => gpio(15 downto 0));
end beh;
