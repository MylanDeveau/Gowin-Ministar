--
--Written by GowinSynthesis
--Product Version "GowinSynthesis V1.9.8.05"
--Tue Jun 14 13:53:03 2022

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.8.05/IDE/ipcore/gowin_empu_gw1ns4/data/gowin_empu.v"
--file1 "\C:/Gowin/Gowin_V1.9.8.05/IDE/ipcore/gowin_empu_gw1ns4/data/gowin_empu_top.v"
`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
ryCze9pA2iwEtOkKiImgNterXuRcyYhATnvfH9r85WuQfXHsn1Z8bp8qXMsEnU+/5IkMIWx3bOr9
Bf7k7UFujFPOdeT93IYhzJBlJaQTx41XHTwNpbRnF3MKThBVbv4U9A3Vtt2tX71RYz9Dnl8tOkbu
5L+W97LPONFVXPzZ7av8fvAuWOg/5M7Mk4Xt/1pnIkVq8FwgerfqjLTLy6Sd5acsoPXvYdzqas5x
jUcxDSuGHxzoAg8yPOL0Lv0aQcJZ1fiPphssE1cBrM3LzrtRWDTdHxbmg6SgMnJAwiQCscR0k/tX
biash7Xf4TRvReB03MnNRLVO8gCiFHXZjimEzw==

`protect encoding=(enctype="base64", line_length=76, bytes=84688)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
h9D3bnSRX3nPUPGVQOewDOtbrpppDpeZV7rKF5/0QGpqxVXxlRSK4oNq8WvuaDMlDYOjr5n87ar0
M4fpfe+2izNDfN1aX82BIpIh9lu6n2MHzgUH5BKxGcR2cjKHM3l4lNf5Gpxe3rSYj1Y2mp3bbm2W
zPy9Z4xBCy+On2dwhwkGdXRmxyX89zYTYZO3/VikYUpyUjRAkysUMZ/gasGgWZdz/rvSfIecBAS5
5G3FcovXyM4y7SRdRxxLsFEAU+mR8a4M1OV8mA2abVj4Pz1Qm577Khftpmmd9+LeTCKCV6UcmiA1
5lqInMXQg/nOC/+8ayd4WQ7UPWWn1n5PPr5FWzmEC+Ax6aW5+LU0Gwmdi79EUtftI1S6lck+Y3Yb
mKbZQ7RW1J15ayGwhcXXaQudzIBKOW/bU2Ny8hYd2LKTCJCLlvJFGnjl54+50X5SnRGtx+h4v1Zq
WonAzNfEDxqo+fb1sHzw3nmxHSiewsInTbsRxXeMpPujjApRfDkXVwZ86Hsq3L8e0koQuWKLr63H
8lT3Yd1RPKmeMCTXPfSWFICfCfGonZspOPAoH4THVv8HA/egKto5x6vi5n044kn49nLCRDias/Lj
ybyfXO9H9qAojL+WSwetENQvRhWTS1LrIIb+d+aBguvjg4/pE2Bh1lBn9B4CD07zELPy2z8ZVUga
oaX2m7Nx1z+LKiJPW+26zXAnzzeYiq9HQF/+NOueKBaBNOlwG27su39CMXm7KwWz9814LSCmX7jd
c17bc/JApuc2pqmX84L0ZJxrG7ckT06n1RRWMwjf5sSvcPdGNamugLEQJyaDBga/lV9TA1yT/2tS
wAJTPOBfYoOQZiDYl56Y2uT6h20jdO+Lr5RJtdjVq42428vE5OZSRkgwqRowAN04bog7oTBp6PWH
led0zKCbeUzXVqiIR9PJAwtXlcy6n54FSSyCQ6K6QWFZsmCTf1ckEU3KwcVTX/D5Ej8m7RC3rx0l
8z8GdZ9EMKwuJlSGcfhPkM4VqPFx7U9OBDNfjbffyVIsbBGjInf4REibiP+tFZiqgNTth2N07QcW
r7Uk/J7+J5xUVp78KPRqfS3LDaqB6FJ9mxS1M+xEHl+MEfPDEzQORZKs9RwDM0uMX9SkXihN8LZI
JmkgrELHMjkusMerjH9lESQ8LaIxq0zTgVpc1bd+dDpOBebLCK2FmhpjfgdBA4IFlcfCDf7JGnX9
QlUmlea9+lU2wBHr+c8pYdeHsKYHXkq645j+EazXZtVtNULLktADuzGP7W7rMToEN51Hw9iCol1m
0d/nB9bZlU1Hz0NDLWbWMglBa3T+c5SVOmgDXF8ylDnozGQok6+Wle9ADMhA7oQKMm6gcwv4o1mq
OyFwZHHqNJbXHNBeKvZi6k946FOBkW1/VsHMuX/YWvJbvJFvAG0m+k6w5xxTCmpURPZHcGVGcAgq
ZkozyP+B2lZchBgD6Z70ucHewjP6R+UwJdfz6whezzL9tvWDwj801ELkCNb/tCbJ/vBcSV2iGLg6
Jbj/whQgE+QQd5KqX0Vt1PB5dv1Wyll49wMVdR0Ejj/dKrhj3XEjazDWiCJGCpH/FI4fns9MP167
slDZtm/bssbm11fMk4rFdUeneABTb8g9l0Gnm15fbCXzR9Q2LFAfveb210/NDvYB1kbIvmrmmSoC
jm3MwFxKqBHH59/5D8VY9bwqKyS0QbpzUuEKWQjmDm0MjZZiBT/hsLNXDirNibdcSLaAkEO186k3
vTtJWTL8nIz/3T7/RNqUUj4dtibU/6uQcKsQtA5th+jT78+W4mlF5AjjQKzsv4iJxpRVbA3RFtGg
FkEKukslPsv2h2Wh/vUo2yUJPU0xt/11mMcOyLoXsljZMe+4bDrD6sLZuUZ647eybzwR3yiRVAsA
rYpPyOH8kv7hM4I3ZF3uupeqBUIgi9EkWX93wskzX261yX9aj5R3klLLHx2MHdMtihCxl/3LHXMM
whTeK35dFEiH4RqtJlFMx/F4l6lzmtTWzEXQQeSfvQXSLHo293QPEW+rsi2kqTbvs3W4Kwn15hgy
T9gysajjpAbwQpcAGhQBMtVBx6dj3vJF1WA3kjpyW8Lq1r5aMeuY+kiOxJfWFhKiBvE8cXLR6Cow
dNfmmmoh7tRT7YCoEATHV48aawPkbD9I4mBs7/2cLEfOPD8vrFYvmrxy+anxBX0rmdMWYRyRV/4c
bn8rOqKX3cNFez/485Iu6eTEP/MTrRinYRR/uLNW8WD7QNpElSc9vEvmUFBT/7e6w5JOnson5JWl
CBD25QLgMF0C9XR7KCVZDV/QoHNEiesK89ej9tni8KjGrsH21c0/6MAaurUkN8KlDBqlRC6h6S5D
CPF2jSoBT2Xz/cpc5n7WAPKygny/HkAT/VoZqQucxo+uRz+BkkvHTLAnvhO/V42fqcO3s2WlGdZJ
5D6TmZGGm4wxdOMHWP39xXhhX9KlUfit8vLoZaPyNhXS9I2x8flLKk82Jj4a6dXWvoGbpcaa8lap
zNHrvh7wFhLenUVn1gjTDtzvWkDp5jj8EfMOLil8R3gakiiBXbsfZKL/ONnAYFO4lpEtkpPcNSik
6vnaT9jbKWFD42fslHlgx8YrPHOumPVl/ONq3hrheByiCsy6ucSuGds9PxvP5Sh/XC5Ro7Ayi0Gh
0cfSXRvJEBuvRKv0qgUAeuT5VctdRzzeFoDo4okQnsrrPsJ3tIwefMlMwDQsPcF0P1l1NdO+Tdki
W3SOz2ecYFlSKn92BTdE7gzE4rSzMs2G+V24fV2DhPmFGqFV1y/+3AtyuBjdOcQHYUPuYzfJjrSM
reuOqXWEjerH58E54M0rbB9yU1dzhh/F5cl2tzZEcGnARpQq4beb+OXio3r/Pft3HYZec3TMMzPB
D+kjQTdbM3d4CX1W5l2hwJhd1MHGyR+cks25fghleZDP8mafCCVYIT0z2sNDrV5N6PFQVLgEv5Fz
nZIt8nvyhvjm5Tl+Z1Vo9sesjfDUpx7hiffvYFXJ6WV6XfCrYQnaCJvVgyHl0HMboFqw+HQpZQDM
fSGZFB5a/X0CqUloNZQAZtUXDpRYriQm5sMb6pfA0Z+wcbNVLGu0S3iS1TsK7brwI2Li/ZziXn2E
KEX5cd7XtkYmB/eNloC1iTNmg0eo/IvWUF7y4hml5c2NCKWadY4gwY0Jh9efDJWk4NsBz+zopX4B
/7kRZruaV9O3I0rTl81uaGq+oql8zp8C6z1BvcUz8rkV1iWgdc0eQ3bD69bumOZkgvL7YEVjo6Mf
MjG247cQThDmjoyjJgXQrUNqkvwLhuqAGLYV0H7F9+Z/ZL6iXxtn317kZQTyQtDo1bN3Q/psoVHj
3jRr/VSGi1N7HV2gA5QKXTlhkfJdLmy4bxjzRVNFTqnhsCGKUF6kaUJmoAtWevz9BuGUcLPYdzD2
1OXN3v2vjMNCTP5nSW5vhatUSx+Q6uIBista2IuKsPskZo7PWVUv6Aso3tVszYxV7QoYSt+IATeK
HgQDEAmUqX2qPw81E3Mw4oyF5GNcDLHdvTCQLJlekVrLdCXvc6RTE2yHlYiXmXC8ofnfehGquTDB
pTCuFkdJRl9YCmBTIRVH8JsN+w3bGpeX9/Hj/5p908x4+f6lMf+qhzGVcq+VjKHbu7yKwPzCVBpX
4fBDScx0X15DtZeYENmVzEfO/n83HyPwgY9QiMrTCg2MmtpXNHXGvjPYeiE4Lky0F5VOW+emKHCw
oMy6sTLMGZkFwsgToAk90Cl7I9q4ky7YQCbrkS/Vg6B+5Fu0QhlZrCI1FjES9o2c94GYaTLHLYr8
Ul8zv9GsCx0gQdHnmSw5r06ObmvP+ZmQQjpp3l+TLgxTObeIQW3ZXJ+0i8KU5DY71NmZixo7evlj
jufhXshfAeT8/xS7WYqsZeFs0dcscMJ6TCJ8IcH9X9+z/TiY+S6MzKFtucQ1Mq+BWOGuwJjZRz5D
5ghkDsPOvEo5xaidEA+hQ3vx2G7SLSIEfLxPrqltzQDvkbIv+v4h0gPYtcGZFaRUfSFb835eH9wt
UZDevg74m7bgA+8fF+XJC9Tee2333IdJyLNdXX4iIFbaqhDlV9W0shstZr1NV9xe7EhyrPnR0C8m
AD8pvO936RQJmtfuOtixoOnRHgnA4B+JGSwLixeDa6Wn++uY3KayYFUWOmSLniX2C5JO56EPN+qT
36/naNt6EurgNROtWuJH2ayRDF3ZmUsJTAxOyIusQvdmXJll3L5wwcQskVoimDNTMm0ACB09NULI
BV0NOME6IP2LRP1L5sBeuokRkDm1ShoE8rOI0Y4+SUZ0FTBzmS7ActVYc8pWXUmxhUJNr6SDS99i
6iXOpcfxUZSY0amutC9ieVbpCGCoW6l8WDzGRkt15niOV7a1Y1XcPMQGBWlzvCCEp8GWykOh9p30
p5/m9AvKK67je5uF1Lb4FKHHKBF8yprhAX2poKIJBKMo7eTGlmH6A3xcGxlLM4RWUMNSMw7cLVxo
wKgyTkPVfXDv0nKaA47iq+SHCliDbsZFCtMI1Ved02sq6DVfFG66YjHELprQzU4jhNcQjGcxN3Ik
8QIuEaAxzi0Q1A7BxG6otol7CxH0tP6CEM1Rh+gxiH2RhJHu2RJgV8aOOIyjTu+nvKxpgcs2gAqM
Vg5N0IdWT5CD7cA1N8233XMwrC8bbb2vEKuZ2zS4NnTqDPxnZkgf/wQHs7YOY+jBBSilbnawVpDZ
5jNKnzVEIZHbxItRc3jOtxCLvAYnjt1wAGV/OnfQ7pM2DdI1BnBTiTKBoybxgh+qbLrLELPJYuSR
+N28W/ZeTUeNNzkFupAzo1Q5SxdkYu2Xf+V0R2i1NqJMKILZlvT40x7l36+cUYq7RR0YauZsvAyE
zgVaWxoIsyI7YW9KbZz5A7zA5en8WQJ5Eo4+LpsgtXMpD7GEd+HBKguUPA65eigPbp/xtwDOkgfP
JVPwbJgwVA71xWce9Gb8ZkC/qYkHDa2jelynuIw4Ae3xv+WZ9IyCc5OAsu8YLwQY28K02UoiV3Zh
tkvIE+JBl7Ry/HQOKEf0K6YODP9xzY+wMROOPeLPkCwPzxKTTdkYzoOXp4WzKCHDa3JxTkitLlGk
hnLxgo2nOtvOy2tIXK8fdnCc4AoMgZiyUL7bjGyQomh4C99wTmusEecU8H05HwZjSZlRAWAXh14X
4sP8xI8Zod7GLBYnz9Hk2N8+IvBOgHFQVDxoKM5bOoyzDTqN7Tpsd0WLAXYxEyRuLgAuqXMesIjN
77hX2ld13FRrwvPvacRZEJwD2+7XTJSvWBDzT9lHieIh+7lW8j41ZSNlpFqSQs7kRBg7yT+Rx359
CU4GIpEwtwUMM8ZeE7NwD2AE/krRHE+Vs29F74xuOcptykR5kIm7VNpf/GwlJeK/jlMbg0MCk2Vj
vcmiBHSZDI19wdJfKG0DXfYpbEQB+6gqEMu3Z7jv78sfMmgkpjEEc0HkwvarVCLTB9JpSVCZKqdx
tGANfDwqgK12kC2kusmn1zpWI8MAkD9Pd7okBepttWd/J4BJP/eVyny1x9OArY4Fi6ZDaiuXINz2
ZzbTRzD/nlCXDZU5E8ZQs6gb8ANljD204zsepIe8Hc7S7mSm6rClcKkGMJE/H9vL8iKBZKCnSf4S
0ubJkwfqbnFA7IA2impdXf+ykdt36HG5jeWIo2PB5fj1LAdlwhaypAogN96QvPrb2lHqE+WpJfHS
BiOBpNWhbABH4pojE30mwMocPujx4pdhP54OWnYf03sG9C7Yex8ThjNBwIFT55FzlWhQDOEP+Lwy
Om54UmEG2LaZuqQ+/7CfK2kDuF3R8AAV807+WChiir5R2/dTtrMrW1hfDyBzdU0HVnDuN6aCNbWW
tIFQk0VhycmHLIzUyLjgnKyrPK8XkWnKcw3DiYaEEeZig4+JrfdcKDefBiytufEjoeZNMoT26s+R
wz36X0xkmOQ1FvOkpXvUZmr/2Qi4FmU7r3FpHeH7Q0DcZWfc9uIEP7ZShliLVcDIX8iUEXrl8woh
2/4buXlFQfgjSZsN7n8+kPb1QxzFLdzlc82u2oArOZSoxjf+PJdXDS7FXh4MeSApBgz6+BzNJYOC
XMeeWQcELnl4pb0l+FE2rVepZcLbFBPTgTiOodQbHYtFrnzB/wtdCpwE8pKgMGAWLAUIvk78WlvF
pdNyEZ6VhYp4aDg0qc+3R6fE3iVdpZvDZZ6uO3hAiPY+1ZXnHjW5H8Cd4lTs6rc7unDSUYdHcBjY
NfafVzfcBRmfRIE0XGoH37hkkNfhTw+zp4dq1XFtsGf4VkSrDlYYxA3ZVCEj0H5+oD5EhdIeUd3Y
TUo7A/KiSuKHxcvXxWZPWAFBYOLKy3p8dYPmHWZkjfj5994mepNAVob8fozQXLVKm+Ak2vqWPxZz
3/DgGMMSFMNT0Kf/lsCl23E9RyEpjm5IJXysg6DO+gVuzNmQQcWlH+v2AxBuK+rXuYMGZTtgCNaz
kdEPyaqUS1kVoL9W5Xs57Mtk3uAil82bN1l9+B14AyNBHirdi7+u0Ze09t6wnH92XGyVBFtpNZ+A
So/A6hnaT2M0tBQnpqYy69QVDRhdSMCtmbq/kYOvxSDFG/QwECI6GWM/eiQ4EEDwZY+U0A7QaNOp
5gLD9Q9TqVgB144EOrQQk9X2j/SdddU1zA7nnn+mv9ySdy7atTKeKZ5Y14AjYpqiDnai/qvz4MA4
B4cq11U9flQUdpj+hljMqvnBDGoC8RcooIY6HwZBmMubBPK5rudLiOyUQgSTl+mgo8qFG2U5WD8y
FjT9SWKjZ1IVYkRvG6gsg90eFFOSdMt03KFTnxQb0Ga58von1p0TqnNMTKvP5fe+6sDcJ8Z5aBDB
sTQDd8KkgwewPbAgngoTLhEenhaaAtnBcGaq4/9A8g3SKvF4JhoSkxJeArL4fWVlXmF7VEbvu5mw
z8DFAajyhRKiJAZzv1DRPARG6JCWoB2ekm4UPKb8+ndOb9Y2hy/w8uN8q/WXSFBic3cDGg9zpjt5
wd8j3JNOdXMUzkoba2U+XSawi0UsJyUZhx3l1EAUp2YpAvl0PcvZhHqqMCaT5FxFP0WLJgRUtU6N
P9uVxh76y8rHl/r6jjaIeFYyOy4wbA0UHGmlq/P7wpS57xopPWeOaXBnOIEn6ry2k61s46enw4vG
fvUmp3DfPZYiXkD1Dba4X1Fl+CTqTvjnEBFf0TNzKuA8ZtoGN079RSZVkVEFGgXNZztrWgd8pRYn
OZcIsVirHxpHtpdLm7LUOrpTjn8vaTWMYNIgkn3Ae6kmYbXLIuWanQawoLQ/JNdb9JAMqsBWvXLe
9y1pV8xvR4HYHIczFGLSj6LaR7bJm1FM1/qUREPcrb8BCiWnhGAYKabgtj6HjPEaFKKVD24dU5qk
ppkFIO7IfBUJGtu9MhEHahcuF4c6d4xeQEf3+yllGxn+0auPVW1rLExa3M88F+/j0cUG0dnP8u8P
FN7aTCYZLbWn/t/ubZ6PkpiVPZaJWZwnxZhNdMXyKoM0/yOdJDO71u58aH1vl3q6UuXo9I5gx9XZ
AnV83G/jAJZEOXBw4hav5h6rzMWW3glrr2jl6bwIk93laXDCQEU/iG6UjN10XoNEplhsIg4KrXF5
bsUy8iQionRnFL4PyqUt8JO5D6iEiugTmyo3canW7o0OIrAj/0DwM40zIIXZdescFxB4bOjDfNzd
L5EtVuys7rIPCU2A4HpE5QJ6OiIAPYnPiMw20lGlgKHTfMDtJ+6Oh+1w+fOk2OIwEV5RPXmfz0Tu
HbgxNaYpVkMuiT1gJDPBkk3/dYLYPINkP7MU6qzm/pzey2kkRS1pcq9d5/87h4ckxCoW1Ps0G9Dh
p5w8LZaj7z20gtlU1/07pJmWSC+y2jMHNANU4Yn2ScjbTRzAvv9z/b3AlfyDQKvHG77vv5aYXII7
2XDSdhJWmuWLM3ZsHk7ER/3p2pNXUbJZxS6AJb9dOn3FkNDGd2ck2S8AJExqc+cMm5jwyL+F01O1
e8pyzjtbf3jmiRBgZ32/ub6kE01USQAnRpoZkWa1MNkzvm63FCOaOI+mrea4lMuE2SJ7mDIQzbFy
t/rQ0/PaKmXbSdeO0aO+qMD/ypjSV+5teeS6IVuUl13riT1qbSYBwaEycaOx3mi/+2yaumYbMUQX
RZ1vIGylrEWm66JpV4VG0LhosOhuiIbGaVVY4xspkezVfv6gU+9/OWphnTVECH2mfiIjGBrLoJHm
f1Np5s9AgKyKVj05bd0rUelSTteSvM1TV19erH0cfJ3fSBpI4PIe3odEWpTv+gV7xA6s3TIriSLY
naeK8CLFrrB+9ljV8SuiTQ3XokVhQBBoVHj+qocs7tQT9oYtMXT0p1BKwKu5PUQp55p8AzuxsjgV
MYE0XcOSXYTYoY8xLvi5ZdhY20Pr+sKit1PPfNhz0xvx7Vud+bRnbijpSwMfVV8PmKzz/+DtwAIV
AhSqriaP8lFtrpej8Y2NDTJB4BSZcGdAi31fc5f+0lAVP5rZ/vccaulNmkpMfnL319kY2haHK+D8
/UW4klTYYDkEEGHIATIcGIcPfttt+ZOEeFn9gHtKIbk2qsS70KCdIqlwuJimp//pJhCEHzZiys3H
mrjPZ7PYVD28zMbTl8TE65tDyMNbyDY2gI5OYFDgKixq9HiVeIHUON9LUvLMCCsmV/pMbmyEaq4g
gXxn1FKxkXQhgLiuZqxgwyQu/64rrClG8zznZMEINgGfAPTWkU9xw87SuqUZiTB11S/Jq8jLmQsy
r4qgJstmoXpFYuMk/3hPx2FBrzfiE/jFMho1onxN1qIX36BPWUwgHYMZaM5Z1Vd7X3BpqmWfjtYL
qWMXM5FbX9II4/7iqwoHIwU+Rmzzh5NQSBgIHiP1f2KiiJ45/eQ935X1wz2vcY0C/hg36J11pVCH
Ls6IfgPGRZVa18EEIJA2CNkRTTjuUbzq2TtaISbyRqKi+nygVMzufHR8WXE9vnTCHILKYv+XZ77E
+QlndH9q4hS9XAzKCb9NOl4nAdikuOF6kXD3QN33VL7yru9IQdGr8SZ46wYndoUcB67pMoWIUh9/
aSn+sTRCtKUZMAWhrcS5mDWk42dID+SJwwkQFE/YERKAueP9IBVKDbEjIA6q0QhL1o5O0WdZ5f6y
i1DuMQv31wkkK/1EdWBiZtdpkhmKZMJfkOrSnvp0zelDMch4Dw5u42MU6zD6UVhbM+vuugAdsOdr
+L3PWifAXNmgcgkcStc7UKe3Bof55gYdMOCegRlcVSQqPkb4LEJA+yl636Uja7gL8UyHD3BW2WIm
b+xdqUisqMd+oRTKF7TYufAHKQyXWLgxF5CXnaYKyYIu5S9WiYQVtGY6homM+24NGm+/VrW7jxEn
y5B5z/6D7rlavuBx7rdwfOZFKBkgxy3eRLuhcCu4KJtdCnFpnagNWJOcGQjatOQpC+NsCn/TGnD+
9BeB3seB5PbVJZNMnmOODRO7M+Nn1NGCTDqhIzjtCKZ+u+F5eRfU5j8oVcT3kayTWFdUMdjLfFqr
vvDa2HntFkUuCKPNV7fLmJa/wMfvOasvRaVZYJ343tavHRG3DqUNxErBNNkVvbL+qossOlLv2hx0
VKyPTxwuQOyZAFqaE3S99Iu+5ammlIpqFTiBlAMjjWk22/QiY0x6l38Px/74Ki6Qofqw87JxhMrs
/a6b3mFHGqJX9f2ddJGYarEty/PGpRY3IHbe1e5cQbI1MkOMCiwzt4HfkijbdKd21pZoyha0lwYm
u/HENvef51JEjgmcBM2WsJSkHfOgfd+N90YzT4VwUOL0Bvs6YyDYMb8Xo5ICS2tPY8RWzIPBuKKA
4rekIhVleeAah3PH8SbswdfPpqUecSOh5Mw4iOsWPLMiZV22IybpHsTDAhebSfK2kGfBFCqjmGYp
vd6eqnqtAKmgPSQFmOL3FTXveB+mGcTyhZ4yQATD1P+DBxt/SOj18Cs8uauIuWv/a/3bTowPsS+m
Ucbg+9w5JsiHcbMkrqnFYHOrdlB4jU6VX2fDA9fUCr9GggeY+NpaZR7hkQvKnwEDSePsvYcUTpvU
isIMiI6MAoSpzjKYqYwp1qv/SklRnEq3GzMM7whSMAMVYOfLjBqjl/2Ct5A7+aRJOwpkPKfPYs4e
SwwFUQu7L2VYNaFYMn5clTOxwo+hffzM4GgI5AIVKb+GU0PyKp9D8Lzw+jZ0FStg4HnW+9Cs4ykD
hcwDTDc/evQSPqHJBHBikaFMcdOjER17idHkGXCl3cjZQ84bzanQilLY6k7D/a/So2VFmWVseh7j
kvxcidyP4dbO2KuWUoUKsM79USVoFmqujIQja9RFRpHMrsvQqdi+dqUTWcrQfyOIYcSzNe/AEkgf
8q8WvelRmIw1w4gqCOI+safRfGOjdDY+MgsQseyWXv36owApEIwHSV6YpuzGInAG3cuxiMyMzlYG
ZyGDZ54t+dMHrD27v/KkqHZiGlzRFPhc6X/6BO5bEeTpNl1yYNLb1+jyj0ZTItJPUgOC8w0n8Zat
c12piKJKUcUM4tX+AV/Il9I6vY4JKwmch3p9h+grRwCKPjHBzZPl34YCqfO20ryyOzTHzFgYCeMI
dH4NmUuaT4HlD8R9emUTR3KRnmtmMVAkfe95d5HMD+6EZsl+frn4J6pUGFPSsXo73PgjrOwe6j6b
Ih8KZ+Gyxon2JyCecUdm1khm5obefd8+nAK0X2QIXe3VZofHinb60DCJe1Wa4Trd8lSs2/rDJxXE
E52OP3nQzZFMpaDEqPHX64tqzGP4k0biFnWvRkjRaXath+ZMFUtNTQMyEI6P9ElLQb41gbjqOlGg
iEQ9zvDXgJ3yJ4aHv5oy+TRur3rWrZ1cNSm6BdrbKtMZZVaqUMK0K8VRcm/HrwERfJ6kCgzybgpG
D6MTVAuTbb6SjZXW9uoG2oC0+NEUNOLuwsuD/DHxlIJafcRiCr5is9aNLNk8Vie/hWJC9SkSdXLh
n0YG53h5uOUHImpm7sxdUNswBI6PCVnpz/VUR9dOOT9TYhtr5R+pfFZGvBfYyegTMPzVFxiofwpm
uEgIT/F8JRQLsrSIJrjTWyDTu3ZzC00f4z1CCl3/zSYnxy/05lUwUe3AGbb6y6W8+6HlH9v3jq3G
YJWH/iguC0c+DPCGekZHhC6b5sX5il1gjAhKC/QUpcDXNdUHWEzj0Np7eHGKltWvhCLhel7x+IiU
MaLa0KzPwrgUpmZlmSQ5pK4VxDCuuzY4VHOMpnaLc5VKOwJhF/9GcPVSPl6q2z4crZ8HgW/pWdY3
TACVnMNM8RxHh0k98MLt0VyzbaRTZ9sYlV4Olkdrgb6QLYY2WZVRrRTwdjHygucB3Fw+5Qbx7BLI
FASkCZ6nWqrL3Wj3uVQ/uo0jWdtNaFHMOF7GvFNA56iBunjxj9lhC6REJgJ6BohG5WFgDF3a3tIA
UsBdXvPRUv7nIItniUrvBdtNronBs1nRBuWaCg71pCC8+JRMccSknlfbKwV6kroNno6SYy6SipKw
mv/5uhRA+Bu3OvlWJtIrU/5QCy9xaryBAlggbeaGYV7a6JGR6dVMO9QEYXegJHo8C8lXrpsjIaK6
3ZcCGsXe5YXHxRNfQuMzb+gxb9dSvqIPxSroiqd677uJBuyld6lCiarZ/Va+xOvRh5R2CZY6SOdH
oS60UufLV+R3qfs/rClfYqNojEos50IwqtWAyfTtAdRETaot/Nps7AIUSPYaxFA5/0Nn6kxogb69
Ca31mPhP8joGIE0GB8uPHum55DQ6iJOt/9Khx+3jm30VOL3FJMzuep7xnAe9Nu68wEURxE974Tzx
qWJpf98CVplA9gKUXQd4RwUYwfNEfHqVYS2cTnSHYLi4gvv4i3Ky47LubbtpPnUAxRuGJ5cy0dhK
3Wm231VeFF8grPkrcTqfcOLYEaN1zcy7oK+tvElJwzuerbvE1jmwuPMZipDMN2ev3Y7/Fc0E2CV7
j2ww6WaRCn9CnYvQi0HdzBYq8xYqWXioyLq7rg9jFx/SyOAT4rLWjz2LEKWle9/E3JZBWcyDpZhX
Lx+L6EtESDuC1l6wXFQvHZeJAjqMU27LtjJAaUW0IbuuxfhjXfVEWsBKbjvmnbp55Vp6ArgyofO7
6grDxlp0nYQ8v/G+09M3cBdua1d2svMjZFAHwfLz8EDM/y2YLpW+jehOBHpeSemOSEYWbsucm7Dq
Q1V7edZtaPWNvx0d1WvLtKaXRxRKn9ueDeHbwOOWcdDaMJv2Ue95IPoyT+qlnuyIpQ4wve0740Fx
OP/+RgLjxpva8ZfEFgtDthD6RGTlLxHX7qwMOVXvCjrRl4ax/hAINMRt6uDkn0GcLFCTFXBiYLhp
rrw3GX8UVVtEjEkYG2MxeMqrmqEdqjLZ4ed/f4hr3HQEwkUKWzq4JnOVfsBYfPX4MQKCT9t2gf2b
pRTxj8rcNusQtbuFA9qpIb9vXa3WmxMoCvGKjmjwfjRSoSEhFmedfA1sh/ZyY5RfbjkDYg0B3Wjq
13QYS5QbIGE4DCtvVVMsP17cF9GVQ0Ud+N0B4ud3nIaeuwOyBKculZsbW6VE79OlzZdG6p+EkiTw
wgHrWFEg9r34T7cs/kFfWzFb8vSy/4up2xuy2UuM9hIT9+54XvGmEU/3E/ANY7mHMmH8T2fGFxF8
B9XYZiTNV8Zg0xP8mbS1LxMb7mOR1O5jUFWqv1hOZ38bfLtekd9eh7OyO2Nx6UG1h9Df+oBbfhob
lE/ZImEEkikJtU+LD6rrE2tfvpvYGI2P0rducMxKgjBdlz8F/0SSzmO+Cvo1azxDjs33Z9pyLSPV
vlttE0JapWKTZHhsC7uac9IdbdcrUgmmhKPVq94yiu0/sebHhllk/j16tnurl07Bl6swC4RgCbOi
dbCyEySs6JOwHOh8jVdIWgtBUZi3Mo0TVckS72OlJTebBe639RkUzWF4bgP+XOPu8Uzg9wya6Oyt
qpQklz168RDCwf556HLVShGf/22itZnANG/p2k6IRn1lxzHVkRajrFbtL3ePlVVFC+5W2b+umHC4
p9HAhXFPLueWme1R5a9PoUvz6mSMsj5Ny5h+WqiAcsjnU8oMtGg/nURX/yIxIXqCSqL/fFkL32Iu
Foqs98kHmId5zajD+zafGQCtaSagK3eJ9+VkoLvY1Rm/53mahL9qhq3Y8rXKRvQben5vlRNEdLGj
+8aqI3vkUr6sE4R5nNjxPlE7Hif3ZvXoX/FI1tVrmyDe8aOYROavweGlGjU7hh/ncnI3IO9qbkt0
qEGTtp1uZ73NTh8WTJ+OTiN3EeoBOGSY3EvNVRYqCL4rhcwrNIEgjAkuwq6cWuKmXOjGOLvB+g2C
fuLhG5sKyz+8XvML42UUr/iA+rLJcz8BuIIU6WfJ1j8GJmJxVJMG5eBnPRYVCq1+X0KliFuDi0fm
NqdtDbuvUtwYG+ip5+2JicVE2+h54Mo17V/l/UBqEJJseBKT8A8bC6jfxHMPL8p5Pa10ARN/tp31
w5CgYrj3SbrPcNpdGxU7y1DQNfifpClYX3pgW1S0u+prKa7WV2nzkhq4e467asVZkBpCKP1Wb7Jm
P1I62HSHalw3cCewSPhqISK5FSpfbNCv65dMEbRkGUvjEoh+bhrc74JdT+3rK15tK2UlmanfA3H7
UByWls/bAaq0z1kho6toNyuj3UQ5qHDqJ476mvFFx5Y6mjuk5EB7+yU9tgAiNh6sj1kHUksWhAGq
T8PfibX9F9dZqvHDusKT629i3bb5lLnlNfyAHYUPt0Mc0JY5I418/iTUthehU2CkrSLAgVi089C4
LyqizYogrhAZD6PU2/MAs+XORXo7iEE6sViQiN/DtFhGDeiooGtlRK1TuhaIORnhUxU9botTlCvM
MND5qLe5qGdbZgH45fRauF26E0jKJ1TNgjTuwuGtS/F7X1QDRzHHbSFbUueej/ogfMpXiP9gdlGP
ItMrkMCRGyfd6+Mv1MXxlO0MNGN+8wEkvcfz5+0bLjbhku6TjeyzhthajrAhgvaNQTzAwBr8Vg48
7qcin5FV5K5TRR/jC6O6/IVJ569H84J9/YLB7ZR4R/oiYzGsB2+wCK6I78VPIiEcfNdIy0ZGDuX1
LDDduJqYLFZO/r9tI8aroyDccAkFxfh0l9bwj8qWq0rX+CmlXWF2Jnbau863+HxmMljjP6rBe7lS
5dohwY7V0w1yVZCUGe2gUvZ//NFTBV+Y3M4j6/N3u4dhZSMZnslCBzTkWxZwWxM3Nd6KVpdt/lQB
ShMK9hRuAH3znrJCjyffc6XRa3dz7qsknxs6cJ3VgD0+Bv/UYMKMUD8LlAOOAF0gQQIsVy6B3LUb
A5IZJrwy1gic5kDayFqMtPySZbnd1iqWC2sXMhZFUv5b+wC3/7SGJrDDiz3XfZoGIyqJw2S6Di2s
khQTCZfQyazhS7Fz9zaYcnL8AirStTqNR7tcjG5ook3hF8fo5HgzRgj9CCwGYIUqO1s99pRLOaJi
IlGgDXjVNoGqalTKPkgkT+we1/MCATVBc5X0BTaccFGxddduYiCGGtaX5wlGB0TVsk8WqF1ZuAri
ty3bJTs6b9I5S/12u9MQlwtt+SVinmxjK+Itl2Yi0XdDtmVWktJKisBOHUJ87X2UDEjyuMxNRno/
LxkD9rIKd+JnpNuSgcZ9EqGxbzsh0K48vrXUbl5Oe9SdZH/9+0Dm/ID7bHZ3MZ1pd65e5WXFThhR
EZFo1B8OKv/MWrqRKUQZQ1/okQUgFI0RK347JPVY1x2cGhMTNW0r4O40kNcZMXAqtBhOv3ivGBIP
57fLxHb8NWfDvlLHuTbqxmnfbdWn2BHI9eIy4z6B8nYGVuj+Q7q+ZC9HSSLhepEqDeS6ZRuwPs/3
kRirvCxbdBGmtp7qcPeFmUJdHPIpdDstzJoZsA8a+vjOOQ1xK7wG/Jx+z9odDs4Eu12F5nw43G0M
ArUOMNzM46yKs0YLpb4shJSBFQZ2IhviyIC+ba9IP8/X1JEOy71f2UF9O8Qd4uYSeVInp4tZch+o
PY9gRfdOmhNSUcF8nOlwFlrefjQvO8A834frn9hfYySV/DrQsXNVUuH+a6IJcM8dILnuN6s6gSg6
iSDD9T5NnGODBgoimv02RG0PJ+Mg/ixrABpdzc9ZvI498BROvm21dNAllo+gWj5GwPtAuLDf/BjJ
A1utenrlovmXV/cyXb67d0OLZg/sLEyYEHArG8R5KFUlrUHUML4SRkgMRElZ+V1jsJUhCdz5Gp96
zubO9sMWkjzPFKLhgZxqRwgFRMivY68YxTRo2pvlHXHoezjiKp4zkd+iOVrAtYJ+fi28MTEuhrvf
ZGNKJjlwng4er/yqVh0ipBUnZMvAZJQkL/Hj+wgr+6valdJFFKS1j6JT4T8ACz3nCtb201mKsD1H
l5cLF1QLungqW6yyERqkprxlbv3h9ajwt3WzFmgvMSgenN/h2sUlB4bKVpQk9W39ftqc+Nkmg31G
EA80pX/ntj0k5H9mymqH/9QX5WvxlGhZVDaabRpoThgFYxqFpwwtaAjO/Q7y+pQMv1ZPbxgNCcQG
kmN/5lCLp/LSnIMMtIX65iTuz97pu8PbKRMGlPNyRWieQBO+hNVUrC0lg1iAPbecPuJaMPEZC/Et
Izh2TrdMkSZ0FASrVuL8X+ssJ9ZvVns7guWrM127EQ8IMq3b/HMutwf/fJhBUDZSHt5C3CNGe+wb
Y7DTWfnC5L0HGVYBKt9/+54kt4WPPbV7vIGXMCeVRWmH/1HcOR0QH1W6fQWUIb4WIDC8ARttNr42
GsBOq8oQBEScWH7wamvIGXTKbwIaK7+woXr0UAhrqIOPr6NEa9rbFEmkwEjS/4chBHo7bkTELMZk
DjE+ZAvtrsyFnQRzqCd/3mAQEnkNvi2qt1xwho02+yrXLKd+QJsey802/Uz36VDug3Khxrb1hOzH
LFfa8svJlW6Voavot+Vkun0pe54DiCqpi87yoSgw5HSuS2XjWMG5ZlSzIj/tHYFrNoAJORrmdU2M
wmkI99N2nPFgr6sdxTUg4d1QBRVZtsNjdXn1+rHXiiVwzDu21mn4YDCtpCdqxZpZ47k8zeBrPPxr
EAcewGnDyS7vlW1cOn7MAZj0ZyiKr4tUAySA0sqiqX4kbiCGTlgl9UJxIF9bOJpruf/mzJ6kGsAl
zMBYqhdkDEwWBHy7r9ZuJBH4xDy25chH6AvK+/nsoYuMCEq06uTr22hwKiPzPJLvsYQjRfl7sGXv
SyrjpgZQXveTUQrxY5Hz5v4/R4Knm9y8WhCd/recONoXzYz/uiLaxqOi+/vss4EznYYqAWQBoG8+
Gzbyyi4FMk+XDYocLJ8Sh/pWvooZeks+QUf4O20E32ODGoXlJMWGj36/yGqYn2cIm7RTPRrC/g8R
rsHmRWINtAqh9IEaAa+uHCRwFm4IR7MMiEH4BMfA1VOzACoTjfjUlOxfIU9FHDzENIJd4K1Ndkc9
8YjQdwEvx1CAIYmWTCyV/0rbPB7SYx4oHNPeTu00uJTqo0MC0omHRk/LbtLXjP3eFtdSUqvHRa3C
O6cAT4PVvONfIyJVTmXkNDSdAE88ttnmsmcP+W0Or8qSRtDCS1koU92Nuitk5JVRGTaA2MRvHO8g
LPccVGylaaIYYjzkyy9Q0c96qlXtLqwi1txXUxTbMpZrLcvP0BqWUJT+Zu0K/lVEmbmIqT4L0lMY
NzEXJkaFWKVtA9tvu/ZqWSbHycIWMb2DifeA1s/g/wmwbmeGMFuVG+XXMKdRq07ReSYSicAiU8cV
Ut9Lm/DgrAo5drZRoe0KV1d0veRYtaUyKMVK2KdUeES08LEvn4Z7wO+Uo4GwAG9jvbmDW+JRLpxu
9PgSUGKkFX8BJ91Nt43nQ1mna9Fwqd+7Vtu/jRlJhkZPXTsaw2OjT0qeFNsXZkg+wkz29ukrdOwR
AywJn3bzqvg+4rLCCsN/G3HEbwhlrDjAX0UVgnTjVY7jK0VBM9gAGrx/rPf+ggDKX9DwVJlo53CL
nmRNE/nIur8DWptKrTSkOzztr/hH5+wAQsqRgkHIyPEwhDePZmRBpO8TdjhTTnzYEodeelPSHzPm
uAH8+qfrEHxgKpSATYpVaP4gS/C+kHlBb8NXGREuGzKdt3JuA2FdYP980fuztBxxfHydtt26Li6a
r7T6r5VjG1uUIwMxcFe32ZpWWuy4HJX2mwZPKVgFtjVoa/iVkqDt3u1MgF5yvJSW3fjFEses/EQd
gA4a/UPSQ9Jqk+mzneawD4SV1kFjdIvFZWyzG1ecEv8g1XoV7P0otZeB552Rwr6i1RRNTIAj2Gcz
7Ho+rVzhY2bX01wdiAFFqSXeKV7fKsCcHrs+Oq4SL7pAKpTutNO3PUdECF1yJ+5IznCD480iXVKz
L4MRt2lSV4FZyyKTU7N1BWAB5mMD6yGoXAwo9NBS+KZfuZnQRHqvCQvIkoAotEymywwd/hvUKbLy
QhuLQnPySZN3rib1LJjAc2BdK1L5/t3HL0Jlyv99I0DS9cYCkel6rVs6PBnFrxY5Zn/hHzZRhaTq
v9JBJ+m+x3638l9DmPUH7DpPtVgL57ixEAVEWxH3cauJ+f293IUIyKB5lCcZlPatxTg69Bb7QOUS
ulxuiSBV9o/vJpCAgtJLDDnnaqPh9uqX0Il3yFDlILM6948+AAKul7Q+GUmxmLEwEhpPjo9kRtaH
hUkHrEuA/czU77xfB3GtN5BKpBcxll9Ls2852UbM4hwi/XTnoKDlQoP/olhznK94837LuZJ8L4Hu
K/dIhKHVpdqUhYSwJCxqF7m+mmV2sngskcqYmDd3GcU4fhn8HOAJSmYbaD6FsE9Ovp6wAS71Lsmb
gcyCCNPsM+6BdT+yRK1l7Pqj3pWawSqROSy6GLaRm+3KiSpjyknrkJkOWx+b3Q6b4FvKYKNUj3k0
Ncdvhrh2Q5mV5srpya1PsMnNOC5X1Z6x4E1oWGAAurk5IzM43IZvIrzRHtrg+4NoSh4rNfuFXHfN
gWf8RQ6NEfo/xj3EOvRhD/0kbFu/7ifeOlLWHbvGs8+5SWtrCnlm1BjWatNHqgWYHAptc7xJGr2P
Fu3oTie2Lai0UsaL0c4sPSORxhdEKKJVmGn3TemTVc5l7QPO0Ut7R7msBQ02YBa/97XluHvHrcBg
7q6cTWqQF0kz98Zw5/PYj6FZ4kT/z3/+WotNSvH3UTO5pkE/er6unOBeNARkflAmvKGRjw7ehcKD
M8wmdeVqkezVF4XHzQghZASzMYW7Mi9pWs5GVO6OlKtcfKQkLcBhMXR92DvOv0187E9VZSzU/VS/
trT46YBOtALEAT1N6tIGR3Dv1h6zHRy65LU0yIKsxg5f/FGqUwPvKPmWjmfRtkQ3NUVFEJZAWOMm
l32HN7hj3qFSUYlR8PXfq5AFpDJ8GeTfLEEyISLXzbGVzP+augAj0pF1U5AbI3/2RbQ6sASjsROu
cyUjq38oRO1jCG+MYYUosD8nZTfGu+PI9fXXqXMkud2jaY221VP86aXlQ6TJ5MwqQfZrW0IzyBLM
cOR6zj5BHEt/3EQ5TtVeya/wtS4ty6hM0UE2WRIMKowTHw+YdX3vk992xTJ9Uij1VXdmRy/Dovo/
QHDC3tnefDdziBRSL2Mvs4Wr+B0YNCbX6mfZhs3GfikGgn2SX9j4qByDZwaGXSs92JRl2tXxC4pY
Ahza1c5yGiYnatJuQIYc/zhPWumVsBYv8/fg2K9kQF2dPlFC+tBaL0ZTEi7Va0HHgQOoJS9IxCaE
97o+6AmI1ewRRuvzTs4kKkcsudfODzGIqrFMbDBW0W2Lhitczu5XoeXKaFby9wgDq8j3HwY2Lfjx
b4keK/3EDVK26iVwFZ6KBtZ8QRX3k/LXSqSvES0+onOEDRetdLPND+Z0GhWxREQsC1x5uwe0Q/nQ
lN7dA4ELuKjRFUZsX8Iw+eec9K9qcUrf3B35N74oDsfnY6NpA7OwozbsYNJHNRIyJfnstsgwGYaX
KnrrtbNbuxA3Ibp0xq4/YOR3XrLE9WS9gsXzepUul0QXAqyQpQpxs7qS8r5Nlg1UBQaYtXtXHgDN
/V6CFc2R9D6z4HvD46B4DJwlrDd9QeB5TRJBQ8IzCCkGxxyQGcLg9BI25AouKAJVTN4+BDSHJR0C
/E2WuYsRQ5AB660OKLN5PWUzg8MrWcSJc1S2cg07b932dSHE4N7H78mKYG0tnc+Tk/dM6DD9kgUm
OTAFjfYBAiMl9/28w66iiv5XKcPZSeS0INTsfkulpAm9OwQEdvN5tJG0lv0Wm+SQXXLZ8YEMFZQg
kxjxPeWHQxlU6orVdHBRnT5Prhu9OiR1lhGnony2X3vGYZu9nkrV2vshN6vpu7a23uQRAZ/vZigb
5rmECKBdh7f8ZXl6GlP0UxDI6ktJG4ITz2eTlqYmOhVSOPp1jhekHaPUsEKRIhVJpdBzce1rlA6Q
15WCC4tZatxfg6dT5WJ5GwOH5I0K/DNgJgvIibLUdHyB2cZdVkeiG3AY4xbyQtWIofhhzatMFKU8
wKaq97s4ClM9VNP9G5YPIiV7kjq18beXJzz1ssJKwx7jaTPWWBbxA7L8NkNmMsxXkes8YBzdvB0z
irMfgbcExkbh6Q+0qGgYua/X7R3oTG+wWVbLzSb02GbxFGogLJ5I1CWTyZMU36JPJXtXLH1hbdSZ
NqBUO/C7OPrP4jXjaZJxTerL7N+VCidji4LfzfEXHWGH0QpCdgbBl3182B9OYYDyk/5UOoSEt++S
0WgtX+xl5AqU09l3H1q3VuLb/DK43g5ZhrPIdD5FRlk1RTAY53lZF1tFlBiK1p7STjQxv3Gd3Cb8
BUbJMwCC8b1UTe0XYDFZc5Vn1tC2y/2ImPeGD8DWKHg8P/aMkk9RNfxfRat+XVAbKeNeZ+4o0Djm
3Tmr5nf6v7DteJlg3h1c0YTqin2WTNX1ThSfNK/50jTOU+ciV/7Q2WOZXOwpdsp0eVwKMxYW4Y8p
yKFXA0nhLdElsY1Xaqu8lxwL24s9elKr4SeL+GX1X9T7bXOQJbiyjxrQWePEWXnI0nw5c3uba7J6
+Dfr4V7mshR9eIsdlhvCNdLvtFC/kiYlxMVj23eDbR8vpXoufFE9RQ+sCyC9vrqCPj6298aHbjjB
q+MEMlbSN8Txogk+wASVkUNoV9SnznUezEHZup6haionO3jXiKzexzqARvvosl9QqhcZ/D4lKgqM
Q7lPuRkud0GUZLh2ytjj5lMtqEr8IZOyveYfMirBRrl2VH0AR+cEd9MzZGDTeQW18JFQ/Li2MtZZ
Q+8UFIZqx2U4/3vJekE8IClyfKy9OfwisFkTIq36J8gNCNmwyBvG1+8Q0rJnKNoBPmnyeMnH/jxq
BDAV89oNw8oJYRoyYWgCLikB4vAhATOwACLia4PoCfQIVWRRk8qZYDhmvhs6WeRIH15XqwW2qzi0
AEakIW0F8/9RCdDjFbZ82YS/vEKGwEK/W2x7qEMAQYW4oQZw3+wM17S0b7M8gDMy0OSIiqY1Qm99
FfWDfp48W0uu9gcf/07aPx96ZOFpPFJ0e6TMP1jwH569fyWNT6zCH56sDHc9pUpg++GXjjC/haao
Ip1BpJASMC+tLdZtE37lvjJde6EngeOqDJzIir0hBk4FD5Q71gr8fJkEVBbvNQZWTxJxl9btAvfI
trw1hBLCBM78y+xUEhqSTQTeLw9ym/Vo6cnA7Dtj+VgJbMlD2fkbky7NHqKR87fjVxrY/OvqvStD
VEyt6NmP6aHFI4CmbG+9kMSrO5dBMcS2TmgAzyh/jO0aHj4K44zN4Q7y3+WXMFAIQKz+ULTlKrQp
8KjBa1qbGAA1FrwDHp2B3uzYSAht7hSw+IpnyBt7iAVZlejA6ygf+w32qf76o5HBXJK3+XKAbRgK
G72jgmKkVHUIzPs2uIDQH2hH2lrlXR1ftvtRNOgUd3Opeg2rP1gDzHRV13RDzN9p7OSuvVG/0Cjv
diGRXrobqfSrjKdVATvUTerpU6lPVkssvqQrEtbUqWITRrhQYrTqnjrL/hw/pIlMl7meBr0yjVlc
no05nxvhPxG9LAst3fPh4DE6CdDz7Y7VF6+Xw2rzS8Z6Z/IRnV/Cf9uOHcBqQ+aXJqTCZE/lTy/g
Aym3UQRzPt4OOcFDG9CKdBfkP6/902sgR447L5FYmt4QkfluWLXt/V2MNTmUvejPqCajvSgIP9Km
C2McESi9JeMLF1Wyut6ZA1aE25WVRwiNQfdj8j1qXnc9jnKq7ZbijCkTQtuZbWLnYnQSoswvuHsJ
T+/7hFcZIXsyY2Pg7bDm9zOIXw4cpcapt5rKQZI/ZennL30iLtfOeeAmb3dpdDJ/HNeKA2MBx5OW
dIYn31+sYN5vNttt2wBhpaLZAt8yR8ZOkEG0IVuXwt+oQk0JQoRMkvY24F87XeeAfOxszykW1LqP
xILBDKrugCcWbnyqkm/CUckUfJLHRa+vyDuGVBhi+NGngK1qIjROtu6rAdaEzEc5slPTZFqTIj2a
r1zMH8J5RAY+LG815Or/KnZS0O5njUm2U8V9PsIHFm4hBlOMQ0/dvYY32R7G11we4nRNt8zJjSoK
kt1bfh7apmtZ3GxFHEsToTKK41UIrOnIsVSbqFjAIVdvrpMfAx1vltn3hBD0sUpab2oIeRoN5JZD
DYc8kFRUT/B+kqe+RjCyQ1coS2HpTYGf0paJI/2MG2ioAahPOnlc9Y8UhwTpxdV0z/NUN4gok3Hh
vxyAGmD1dIxzHLFq0Kx4onTots7t2+sdXjRpg2qZrcLnGPOuxGw/UDMewW6pmOUkjcHsBNkQ+4gp
qz7bqr9KAODOG8gaRKmXLUPalBDubJko4pQaiqXEz0o/8DWLDWIQizaabYFyxiTc8L9bds0QC5ll
783w5VoOEA4bITPeKOm514IeUj/QnUE4xYVth12BuDjyyw6kAOgA40/0zDYg9wskYMbzzXDXong7
welL4l4E8HyHYR7g+vX1/iMH6lwn6+e3gh+heGs70NX825MtF/9w+OrA4mByZFC0i+VTwFGj5rpZ
Fxp0plRjAh9ARnCk65L5yxuqBPnY4d6vaRA8m3ag9QsABw7JN6q9zy2t8v2SkBVpr5UNgFIr7a9a
prov8Az8InuE/LAh/CFaFxj98vck9MuC9TZOWNvbA3RluZiAAQtifnWWZJYpEsxmtZYw8bAD4lyF
oP4EHiZiI0lhiymnRqjH+3fJchZ+ZcEFUd5qEdQGiIFeem7Osgt4dHZyttgcrXpgruBJqrN94ljb
br8XuojA36bmYp6etvV8TDfEzjlmCMseOfT3fQL3JYT20Ig1IfOfGuLJM/fWqFLB0xDVtXMs1X+3
NqctuQ100KThbUTbEUsSws5UTQPuHXLY38H9MESrBcGy9GDke7K6D8YqB/F/BcAX1GLiGc8xXag9
Ap9jtfecWvSHVHPF77yqULe8TzgLVLbVBSaKOdAqPa8FRkPginBlkWrqMSkKchnK8KBK0sb+6dHK
H83msaIssXrA/cdUWvdM/IMmOhaEvlR1q/eAAY9ZaidH6WZ45wnxOV/yLUgAwmyZiG9MknxjgUQd
dTob1XbGdESK7kaDo6D0OPY7U86izBOrbiNeG8G7lywcErVMFHmxaVZ4zc8igyisozDHgSHF1TQe
UrV+5BvlThj6icNOhWRs4cZIAgp3XTBkHYDf8LOz2IwijTLndebL3XoAk4Vd/ou6dVPjnCAo3hwQ
zUZo4FJY21GdviRJQPXeJYX5SoVHb9d+k1sTTs89KZzbWLITMDoJZKuu1B88Fop5z+XpL6mccnRW
1Py48LD6fBjdkDtEb0qfoQ3ggRoprivnZYJZo/lt7712RBjbmYyOJMO/A+HC+tLDbQJqJa6nWEJz
tBggLu+mWpDGJoQoCP0c0Nyms/gLHNzmQ/aQelf4O5qtmHTDyTykF3ha6W2b/YaU9iHcPzMs0Met
kc9NCTrArWEgTL3P1XyCeOuDVGywY2qiqkSLvA68EBOkwvDDDMXSQ/jwzpop3mr4tIw4GM1QNjwV
I/HL+SswQrrWIu1s3mQ0L1IX6xdl8DOc1+5yCTClcwPkhMZYiepVJluKnd3bl9QewKwQL2MHhRj4
uHeaSdytsePva6nfpgEnzPC1hUqd/+AJdX0oeBRVQDVUK0cd4gN0DhYOQklrr4m/mvvUkJGpji2T
Hw9mP1R6OH7IxKrvhL98ZQJdY9ewZLw0YGB2Agna14hzoFS9vDpz2jfUxKy5YaMIPdaoKdJVOP0N
fWvpS5L6LyvvBahnjCSLUP8M70ppiihlbPj798keOtTbu6c33xt5rA+DesFI3jzIrk8wN2uJteFl
MXNzWlGViyoE6HKcIcYCKQ6izsFc6Nb4U+TvJ2LSog0MmO2r1sCOxqwOrA0phuobF0aPiVmxrKzP
j/kg34L4Ef/caA2bjv7wtW5IrGZY12HqgGI7EE9YiUMvIpFmoFuOU692HUI4ddBEVM33P8eKlaRG
fbkQOmRyNpxRccGP5gLiHbxnERXHG+krQS9PO2ubW+zunaRepp6EmGrOpNwMWGB/bHG/yzQT/jhv
3kJrAGe8Loskx2QxblNftM9O606nwri3vxVjdTS6Zv7Wyy8OlNmS0i+6Ht/ZXTRNxwrYwZLNp1p5
Uye4VRn9jawDuVUC9MDPSYAzDXdj68id3BL1Af0xnYrv0L8HqgYqZvj4eYYvDXnVwpeLGWrU9qQ4
TmCgw0kSX8z0jXsJCr2dLudrHf8cGglEmut4UWgsEQh5/UAd4UWp0R6ZDLJGsDYhtAjn/4kCbBIH
NuEdmNfyAtllHB/LffAEK/oWjZPFjKOiVDP4GKShDSoRffh2tNz2UiZ+W0mbBvmWPv8LBAZ824u+
hfhN9LYUOMJ3bb1T4/fu/dDPE1txhs0MZWJV9qPjS8K/Sd6oom9jC2FTTWRjAJ3FBWsHVqIXBYQA
sikzxIw35yDENsVVjG7tl/upDEAX8Hv4kmP3zUCoTWxhtn3Y+dGXZAwolNHdrzAGK1StCYxDfTEL
SV+xvIF5t6Q4vul1RfQO99kZaP1QczFF7pBTpseGo8Cyljaen7ZSCurOqvmvQqmDdU+hLsxRTtWF
nB3x+PFVsA7eBRYuTr5JoX7fSlsiz1eh22omREKylCKYxw8X3NrgQe+ESa0BpbH2q4uJ7Ie7Fo4o
lkXLUigU1pClmbl0BBTx434xzDg9DKRd+W2W5SCBe1O5ybOD+MMsAtPnqFYlrlF+chPnXMn235x0
dyPl/5nGKHkDuiHp9xOmnqUIeRMHV4wYbRhmFt6hMuEtvJ7EJKCYUkhgsyq7fPr3BaNheIOQi3V7
+UAEd/KVO9qvMqv3ndWF/0+3+sPXWPt26cbVjNQW8xQlzxlT5CCprIlCpPJ9sNXyS2XIUZarlPVL
SAV6v1C0jyAwf4bjFNYQyqHwVs2o5SqA+uXhAqG1ILBwwLt8Dhx1Qu8mZ3+kqTAef+8YoXnsXNyW
Ilbgm3NBTvSemJY0xhazSdn9oMlCCKeBPjH1OC4nDlEBuSFQ8GOPhQYhVdAYdYwU8MINIYcnBQpl
bdblDTCXc+yoRLY+2uI60z9rQiHkKpiuo2m8XdFoYPNgNW+Tw0XVQiw8EeLRM/84U/If6J2SEvKK
UbNX6gRRIb16Z7kAphzQqAXhlcq3ChIinbnrRpDcHw60/hgJk98XrXKLniHdWWToOrhjue87njOL
GWUesyUzikqBouOk8WG/kP+cxo+i0GTTdJWL1SKnycR6Ol/UI4uR+vYkv8CP5zADYavrg9Ksejmy
fy0XlIDGMbKoKrTzJ1SHDjTGbd66xgQqIDia8OmevkgjAWBgV8iojD+i+WAaxTnJxpmzfnAqDLqo
ZF3n1CJLG5+wPx7m29WVJMhfrzJsBxRuyelEuQPnjphB1DKk/2qFSvC85uyozF6skoir/l8w5Gdj
cAtYB8LF9ZVS+9nuSPJfPve+aNhdeM7hNoazX4JVnAxtXqUYnz0P0h6flBTXGL+8NqolAxQi42dt
d/vAlbtCn4SM18Ro2JVSoCzBfAgUECicoaI06FvW79Pv3B8KjbRfQ7gNAx9L0wheA0kMdgJokZyb
Bwtl6dh9i86bXru7vaQRXoobdei+ds1uq0cbDnNdEkotFs/k8D2pZ5E395ASVmhrpRW9er3oZGX4
BmSnKa6usquEsOYrk9KlhaFl409Cv1c32XbqvAST9ysAXJ+JGjIOcobuUvHUt0chiMzLjXpew5DN
5n6X1ENS3/GoMj0xI7m+fdA20X6u8wxjESEb1y4oX9my1QT81cwpkqOVAv119zilKZlEN7R+pU2h
5sYykKXFLe9/ABEtJpBiNvXfTHbid4rdXqONfwUkBilfh0ChbmMMluGfcHcYw/1NvD0IHppfDtZt
bhxExMWxQXaBbU0gXsvjs5Bdabv3h9Kx50adeqtGGdB7r6cnvu4FQDbZ7k8WKgc1vY3KhL/pJmwr
gVs/5Q3sDlDVMH0FV9QoEe455+bKGsMGG80AmeOHXtn8QpomzUqWKvkFaLJcshGT5pTUsx2uoOQB
nMkaDWE/UNFaK4w0IZZ25i17IXeJ4Hx+AjSW3KL6Z7nSNzXNbwKkOwmKn4mZ5EWNS96TbKi8gXfA
e8YYlvZmvarUsOz10Ki7wuLC9tFkjz1RRjs/GdVWTyw0ruVTuklNkGCQMCT84qs4dKpCGPPZqy6N
+rdhl9A08PX9SMSTD1IHZB2zDH3qkuBNJTIfVZbiKnMJavpX2iIfFgJkv6KEi1qkTA5NCkkIy3D4
YuDWIcMzG7T9fxaGOGDX0rbIiDyFYJfyMRYs3h9mFxsukvona18VBnKypAnw/HmCHtF+dgAZlPBH
uiKzVSJPab/ErJ7lV/DIPBArVhk++zs4VnET6JUdNCz2IzFQb3A7TknjQrrmWWQ1kYeuQd16Lnck
5ePRPd6v8gREwE4sCf/OVyqyeBxXidaIaqjo0hm0scL0u2CM9gP1QmXPJeMWi2BKvyr30ciygy/7
o5+qVL9RqwVybda6jhNceKtksvP/UmlS34mzGFsJp8bArxnwVCPbCFk6YTsC3CukFxGELte5pZF7
d1WxuXgZIziUDLCwDziO5kWgyaQXjk16bE6cF/Zww3iuomb7HcFZDlzf/IqBWJp479d3L3+Qv+kD
Ewd1Ba2NOuwgc4cholb3JpV7QPKFH6viko5Gwnn2xdLmnhMx2fmWTByAb/4ka4lDlO56cbOjLWri
FZ/7Bzp8fbmzbSAMNzmC0sDdyku1N/v/36PN/ynKbe0nbgNsX13GGXdbi/XnVJPDuIcsY7n4M0Sz
pmZuJvXhbKJHAHFht8IMCVbPH6w8PLd0xcL+W2LgpB78/Gj+bKntSFzNhVR7PEX0dBLg9TX2LjZ6
nCmcqx52eaidvhiBZYxu+FptSxyWSmPDVG9bCwyK954Cyia8er1ofrpZzXAJUQCh7qYoWwB3rDKM
PNu/yPdLKdWFLOcmUQAzcD/d0+6CYBB+VjGJD7BPBV87wf74YtiSIyb+jTqnDJpXPhuARMIygj+L
XeAOJ/i1Uw7H9vf/P/EHUwCMLCj4JRH8oVpfaUln1bt6J7U1sgq60RruPdmAwgzH2laZ434OCYzf
McqcbZi01DMO8s0H8yUjXNAUVssvdD2TLYpPmXmpZjwnWpxzstzu5UwF9NwJ6MZL23nWiKUcS9jD
J3AfMImMffdGz8w5pGKGpNj/G90TDYPtTo86v7CRtW+VCor9Ne3BX6vH9fBqO48ghevE70th2KNF
OHn0oxshbmrzGrDQnBqzGVjWQ+qNt5K4eX47D5ohILoYerqjHSYtUwXbl6I6PsXcBfDP/8mGmuKs
JwnHRPnZpHfuMB6uPMgKRPDWgKoIOjjjW1he5GDtLd/Kfd/jKz3Qr7jGi32ny4tT/J503VPDtVnq
sGC75opI8bhqinEWb6CW6pSxthJWjqGZMNPFKIHoSxy3/3v5oqQy9H1LNU3O9wUEoAjL+XiGCBFL
MPD6BofFvUaKOEqSGf1yPApQB9OH7aWhFQbzYirIjgisfNgTGhokaTH4R/Ymhw5qYz6psKCauosp
pheSV+t7X4shLLCUanGwNtJgCUbX+rfx1ahasrOLCKr+ou12OYY+eEdOfCHFeoFstKSCVtdpwBuI
s/73+CyoNGPPQ7E6PaODt8E1aZ7E4zuEldMBHwfrimDIwMT5TnvQtss5IUtiO/uKbELeKffRqY1o
xGUVpH6he1n9Aod71SFrjX6jPXXeH2OY8ysWRYCCq5JWOmbR++lyI3uZvENgS/i0kEt9AGAh149v
LiNl8HpMVtcIxFlFddin3oUhLdXzajHzY6ZIhKYQgr0UOD67VqsqAmYamyEJRNlZ57JfPEKiQwFr
YxKrdgdxFLW/eXy13YRLANs8Zk82N03g3ZXtS80x7RPbW0OiGrt5EWDXG8J8FOznExFbH8vzK/ZP
q7seM68NPOEIJMmCZt3D/GEdVKea9j+9pZ4x4zX6kT5T3I4sKmIHAENvi/Hj+ZH92q7c/uUnpdYa
B2DeBVq5aax/+hfujg4/DWj/K31buHySlHPoRv4qzxwgqdGPGy51vXQZcp6Ibt+hzo6g4+2yO0ru
b6sJsaueFgYg9uV9IkBcPYRHHdzSn+ToFnjzfmYu88ObwCkWDqqeyQQMf+W0tqpsn4+QTwdeTXqp
iDSiXgvjdW8yPauK8ebNmwfRcBXdtZ9V34sKx2gDuOe+L0hMF63DmEb0imZUw97Vu1o52yojaNzR
qDhO17Fg2PFs0u+J/aje0k0uwdKOfMj6ERsB7JZvRZh+LbdS2ftZlmhGN/hN6wYiePvWVwNprjZX
Y61tf7ThE+0/cQ4pPLvcdCW3GAdVPMOV0nuBQoDy/kV/HBA2n5WwpNos9dizckp31YAV0BFi8QJS
he33KLA9b7M69LviXF6Fh8Xe6zwDcuxBz/nbzEzdDuP0iupC+w1VGhiIVhvK2YsW3mYSq/DMdsLg
5S5vKt92wzXem84hTOaTbDboQipZaJSAxIgFbvyr6ARISH8MfeFwWOzO+ms7UoJ92LQvz2hqYZSU
3y7V36PPBIUxZ+yr/el2WKOt8ynQtPhokESpfssivtu6uYh94rj3JpkadgFIR3/x08hQws8j+fmn
zsLejY+PJfAZV8Rw/GAENb1jceCb2HTTiVhHxkoDwoKMm8Xjabk/gAUCbI24WfLTafJd530H+ppd
YtW+tnxS/UdwTwupDc1BoI0pDInU593X56oApMgHpGxT6vP0VDvZAPkikZyayDiQX/fOOHka9WRd
wWvHIh/p/6ONNrZWgW2nV7QcgrqtVzEN69gQrulpEESVuccL6D3XaBiA72CkiM4BGKj6yJjinnpB
fmQsNN1jAhRiREVZ8lfMaIfhXc7CGJShVWUe9aijbNwMZrn714XNEqyoWa2sY5Z16WAYoPuZxL/Z
aDUwB1WiPu78uCe0dxRCla076CyQC56o1YVBJcsNkvrbQvh/HejO0mg5lI0upphAG9rw0CFXP1F0
3GWmRZ0f37tM7NEBjtt61hfPniMXEPIJi6qN2Fgtu07qZWNmZuf1RcsLNXdHl2H9AhgAoS65YTQ/
uEk/5CLSyiCCHZoWAUkQ4D3j+85KH0con7m0cSu4XQ4iUM5EYxgYYToeAK6h9XgYY8HQKgt7jLCB
gqlY4J3zpsWe6qKyoC0iPU8wo4NGuvQkZQPtaSxzuA+llyuR6HUPrwlzuoimTdafxwKpyO7wnK9d
rc23j88hcdMM4r+k8zBiD+VYGSJK9aalVrV0zqSWsFrBuHcxk0Cy2SuuF8qs7sfPrMZTnEy737Tp
qZn62Z4RDoEqvrSuEyq/71brYN+8Xm6z59xrHuQCCSCUNAogEB9pd5pTwfLCxh1v6gF4fDn7kUk1
KWKg7etrd/vai2m+CCel2p8lGLJWqGrb8eSo0jEjoPxkFDg/M9jrstLi8busb4z7Nt4QZXVbNNjh
pUt71L0KJttIWKALJKbf6F7B0UrbldspkGxWpiGvLKsusVszrJydo+PFrfX3bAVkM2Oh3GVUvoIj
nRyEbS+j8ErF2s2g0IwwqdwP+1ii45E4MLv/+PNwKOwrExFnE62pc+zvWNHBE8uWSiU4MYFvNqqY
Vrnr9VVMpaoMA6G5GsYm5wK3wwypbKBsgZDXlQ3bLwjZ1w8MoEWNJUZTCUI+8NQzI5UluJc4/qJb
GYvKgW/BNB5iigzLb6+4gTRUko/XeNcPqN0Q30ltQ3I5NOwx2PJ0VbTE9DKLhQTemuGhSDboczSH
8GMZK4J3yvI0cpzBhy0K6auqJNH6SQmH3TQwya1zDbRoE57ZD7FqQBZUH4OLRzvwgw8BNnKod+ub
u8Z5aNJ/6ojps1OmBN82gZTX1Dq+jjIFonGZ5qL8LIMoNgEefUM3aM8DPmIeWKZe/GsiY8BTXP3G
e2bpjClIA+LyfJMmYc9Wb1X//4bFX1yr5hBOfFMy8hFRaO3Lr/S+QxZSc3JBZZzup+V/TH9is/Ca
5xfMvyWqTdLpZwriyGScUgArqAvXw13NvXLApUckmJdC8aG5r8VZwUUHWuHh8v9CUXA/N5n9bn0z
U9XjKmbQ0wuBjJmFMmJzTAqESkMry57I3ybWie/80LXLzVu8eYaZz7KOqFONdZkqY/ae2J4EZGCz
Q3uIAPNAeO9gKaYgvCJJdArIu7DdWKypU09NBU14sxGB+7KUN48w67PQWo31bRsfXHX61QKaB/px
jfWecQYuhAiGaKM7r920FhQWK6xONlFQ7m6Xu+SeU2LMEw+HsE0ZoRo1SDLUbB1diMlEmZa5PIoF
1vY5hwjOlv8J8AR3cDmNnLhqEeeJ5gHdDDJuEO5V5kmmUSMd/pe1H9qzFquKJN0T8YEtNEV6znxI
Zdo6T1TWm9kOuqsTKX2/gWGz95RzuMF4h8WFdhNcoBjde7FHp5Crbe45+aGUaC7j1FqDuFayaZ7J
/5xdTU8nwgm+xQeyvW7igITuL2SntMqSU04ztykE+fXPtNrPeWD/a+28Wf6XtHHGQqgM9OEMLoWi
EGLzK18yl2zrp1c6JfVyGVnuSzvpILdnzNEhVr3gCsERYL/zsqczj+5fZlDQP1qHEpMv0tWqxLFs
4NS3Zuv+bk3B8+nyJ3asj6UaubRivs+z1kiwSgvLrqvnXwQtPJu7X8q7FeJ/4hAUSvmTTjAWDSC3
foBgT5y2IWTp8exXzrX6mLLKYgG5iMOdjPwOF1z3c/w56w7kQ8dV4Hr6L+HKni7AHNHhgPiVuySs
MeaZCtBAP0JpSsX5pwCHMyBMi27+qfXpIQw8NGfZLzdfkTMwN68ZtTysG4V/MAYIvvAD4olNr3de
ONNyya3sOA8Jvve8MAPG2SDUn1IoX3F9S77Se/mA6kcgvOysuvIeI/rMFWenpDSiFLE3SlA5UvMM
7M/tsrb4CufKiBiCG5+uc4/nKVWQadL80eEMPXOoT5oRN29t8bgK4qT82oRS/p++nqXFShwdnCDv
0pIMnAW4VYDICHcPnMixLi9Tk6cpYhKQ35C87if9r2ad29/89g6UkJAQ/80T4I2EjNOuVf85c+zs
uM6aNB5TvKh4Qv6jhJZH/3YZf2acfQdvw0eeQuNMLTy4FCrqaLElQdXsxWJzoweitWOaAA7IiqEL
cjUOPLlQ4VFi5C3PKCAa/p5/Y9XVh14GX3FHkOiwAoSeGmHLExfzbdKPx7elcMxnDIFmG6/8Vw4w
UKOq7ieQgyHA9DJu/dilyvUiWqjWWOIDtjiZ7GwjAtwK5knly2YmngI8DiRe1Oa81ulhtKicLqsO
QfDkaS5uCEAw4Nz/5/+Hhf9D7p7EBNlH2bdIVHdq5RU8K0XL1Z93Vyj5oWl18UgMIAHzVCPPOiGk
Yzw1Kz/5lJJjO/gdxoM2z+dNfkPKmyBvqz1pA9EXVk4tpECZq5gz1kzg3faZymU3mZcWqa0K+SS0
Xevxi9qxWbzcvFmQFOt6a92FKfGdMNUCR0A2JP9iXBBt+TX8ieC8j5GHFufeCrgH1Z5PNRngRyVw
UdbsoIN2d3LFcWeA3Pj2CkWaNPa2tJKJtOOaC5nkuvvJYrzJHT/KhWgCdpsLGBmyG4cMzhtzzX1d
wTbXaLzBS8cZZ5Y94wEqef2fY0A6T3hGYhoYhPj8ghf6aBWEEBSB7wBIJjUUtD+tna/gN6Fbrulh
JzDtJ1tN9cZke/TzFMES8skmBdaen+f7p/gklTOl2tT/X8dq3FijSmtxv34E06vconJoRZjryFoh
nnATlhKnr7Yr+KmraWit2Izq6rus9EgJO/uFjwgLMVpk59/djzwNK86Kmd2dko1jBpzwThQjleXg
aNhQMUz/Omyqg7fDzMkNoVQZ0k9LS9s0XIgbRLfnyju7MMgQbMYg+jjFPUanfMbPH+eo6HVRVrwU
jbSSpc/FVUCvcBwLTTAqjtXRDym0aIPH/MgSPhb666/P/ahxB1I6dNHkutwzXvxURvkUB2k35k9L
bU7dZHRHgbeOnMH9K3kfBptwNkQENfF20y1EdShCMu6B8+zm5C5YpJIDuTxHYEbtyGRdVFD/A9B5
fIBDPbe2OuCKWyDuD4QsqqTcEzt0l4hDTkHQR0ZYCSWbvtvCyiq+/jmbXvX6ewl+lRus5/E6rNd7
fEEdkNxc+4HQ63Y4S0KVV7F76RJVmrTY7iJQI3Sbt7ggnzrc2ltLDHSiE5XdaagSVZOiha7a2z86
U+PB1Cexpoe4E9oK7bOoGTz7+f3u+MyRcBiHB+FK6F5l7nCZ6HpSy6AsSOdaJjfyXH+Bs0unywhK
hgqfpX6ABiaL5ffrIuA6nOw9+CWLqL7G2a7sbhpJIcVYCnDYZrvpvXzvWxzwOdXvIO3TSHeZtQRn
9qKI+dMx+vo6GqXH3dngQumQiQhdRHe1yrzCCZvebrgtIplwgeFunGH1pmi0lpx77tq21gc/8UBL
LxRCGhfPk++kS14uWSzBvpz6oKvsj6dg0sZ5dUTY+KEo2h7R6yFxCEreEg3BCtUiUlNz0eoJN0Jv
8V8x99OlU1Q2kW0+V6bCLf6GRk1tyPgr1Xo2wF+dysTkssRVDmGqARhV5uQUrL7aHxYLIf/pi8jB
lEQcaMbXlxJ/Sq1kaQYmeXlJGKD1jum6/1xyrnpMbYU4gkTfwjt5deQi3HB7fQjCP95NVPL2b42q
ovo31lpAt7jFRxB5MeoKyITm1ZAXhk6x19NBxeSUvOtL9cj79fYJ3kZluzDhk4yW/au4JDycqVVf
6dGmOJa9NAUtsnVenegUUIKqE/ZVwBO7bB26FzQQw2QdtML8irFS0/Y/0q2Wa8+YHMR+181EF7fw
S9robQevPHlyUvklTUx5rDZukARX8Ln57wRzKfPjhtP+MBh41rKUVdBG590PrCRe/xIijF627hoA
F1R7Bm/MM9mxuE3Icy9j4JiKTEVXhOj8gHExXKlmP1bDEMA+rMxqwNchYhMtpBclo2Q8rD39BwpK
/Z27AuuJ6uTA6bVCCMVCxihMMMg+hKIhnMuMbZ8idsvI9+mp2ZydpjrhTimWEWK9c6mI/m/Qxjmf
F3WIuFLFLDWLczjL2keX8C1KIMJ9OTsP+aEuZC3TBfk6Hbo+Ksl2MIav+tzVfRa/HXsy/3K3Un0x
Hs+U37eG0yJYA+s5zNw9p4jS6U4FQlb2O8gm1Lp21Y+uyZm2qv49OzFUtUcfddZRf/Bk5u4Dg1ym
ImI3end/sl24yv0locxNeiEYP+171EEhb75wA8WIQzZvLdi1yE6+MVGV22qj7DXfJRQlEDX3yhAz
XklGoqxWONRCw4hdIzZD1J5xLY7RJjBoYlL6RbRfDgKxPDgJaxvwYeSglbINdw0cao8nFX6pZCBF
fD0JNRr7OA0nz1+v3W/t9il9a0rK7UFLpRbM2LRCgEWGx9sGLokaB9qAsEf2IKGmiWsGCRPJlkxU
EY8vsbaBLIwwuis3IE+X6ewmnGIsmxtoujRNVPJZ/r4xmsNVNc3CQAiCyV/tQyFxIZY81rO+Pl+d
TSAOwHqKJZFp3YbmeF4XCmDf+xb/fsoBfC2wSONPtO5QNk/J1COt4y8WcAR+Ir7Qf80ujSPpzGgR
ZuqGLv7Dvg85O8XXMJUmLBguvDu9umYGRnTJeDfIPqRVTOYKAowEqu2ZvtKe2Hw9JDEckhPH2mwC
KuoYrMQNbYJkFQkXi9V2gHhaMZD2ZD5hVWlFpJEhdD1Pq+keUkq6ME0I9J1dasdbcnGNta6E2jYI
UlMEptlXIL03ZVWQyMbVVjJyliwVMY0S4YP02qRbsPqnlplTHl8CD+s9pcEwfsoBp13CRAkFbtrg
tPv6TYV4LKpXRpgo56vWx/u+80X8RooZSxDKKd1oyvfUwbDNM5PM2HMth2pS+rhF7MPZQeSGg3kk
SgKqnxoTVGHQmmqCpxzLu6gShEJuPLvurj86Vtukj3bkH5v1ga97woCeJr93NNr2FqUl45TIyN2A
pOGilfOXBdDTFxc8rRXK7YhgCM59RilKXkuSJWL1yyL4krr69yXHLG/wTJO9Z6r8BPQyukUz5mSO
UpOSS/QBu4ToKnfsUaSwvYvYnntvxVqcu7bUoutbipZFlmobCsPa9HERvgxlMc5V0b7B9UR2lzXA
reQdbf+AMlQdV4JiYKMqaMWorvbY2rNSXACNh4nvtM1VBb3HF9S/nIthWvFILtNjETKVkHZ9aNHw
hO5kba2HvhnM/kvE/3OUH6QP6c9dgoXQeT28ymUiie+fzblNcdV1nyqFTRqtrhlBjMXmFzvBGqVX
fOolpKdsl+tyQxUKSTklxQp+uNZ3BiloBbiaZFjFok57tG7ykmeNCt2Kfcw5loF9Uq931B+LKyNu
2LEd+2KhNEegBoxhw4iPwCVFuQ9qtIS2o7s7rIpKq5P+W+TDhP9WbY1/8JRZ+WawXwVbWKKrNqQC
HQ6GFi+iHNCj94ifaw7PVtC1nXEhG3ETuI9OoVD9VUAHKmz8Og+s56zZhe8R9sfqi07CVyMOVXFl
tzATXD7/k9cvhgtbNNSqD+i1MGRBNXAC9On3Um7C1n+uYAugLPxg1eRErjmTNe0EviD7V3k7l16b
QrZhRkP5w8fLd7cMdaObeS3z4K491OpRiTNipomp3DOtXdnjK0jeVVVpbrxsmK4QjQ6Y/tE4LKMh
HjdPiwWGOmvCTFq5ovyPEBdSzMnAX/KTehRvxcz4x0dKeEb/iXCJHNifsUPHv/EH5gQZ32UwtA92
yVw2V9zafmCjdF8uMJVB1i4hsWT3dvg8/ANmnP8VQ7A7hUND1lPBy7ZS0XQln67a6lvwGHhGHyq6
YRc1buiYnJ580UfYtbl+mjcTdy/xH3G2CFwkD1dNyLFMf9Pserv3nCCpTpOD6yQrsMUZ5HsDThLW
8Xz3mWNlCxmjvfEyeUomXgF9cw+JlahkxjsZXonTSlMfRfwRa3PtJ1f1g98YXM4umOW0su/YGGp/
AXmbnErv0g2VbhotvLZ24hXghXTN//8PWMx9aL+C6dVUgwAMuSV0At9iTSzW4GI1cF9FbAFufLfJ
c60AjpIPinluFVA0aZ4G4GbEky4ZxtIaicvTxPg6tvG7L/2WePLaejK5x3z81dfQuyb3KLKTFkYd
eytpAgaC2kPPnvlo/iplZxfVeBkKvaCdvufbHbPo3GPdZ14sQKHaoKR4nEysWo3FfqCK+vPJRYV1
6OOAM5YBXuBlnS26ka6PYjQiYQ9/tqx+7MZCUgFgdIWDLVbWJunaNXDuB9e9SOX+7QQ9xkbBtZBT
SAjdU63MwcEylmd2+UJ5HPAOM6Zl6aA/p4g9GAg46MQD4jEMdSbryEroRhokbNMDQbQmWmDIt3d6
MvqLF3+G0YlTYeZpBxAvIHQSqiuESJkpTgtyRLGH3zq/LNpJJSd6qePp+xjw82bVAygMy3FfA3WN
SXsIPhq2jYditKiWpcUHMzteNZZhy3wNxoh1dEfSqWkkpOgkazdD/0s9H4nEzw6lPLLRgvwyY41r
eOrAWBHkSC9Y+l2wFYmc3hJGDI7whrhM8uSbAp94KX5AmZ3Ur/T/mZwR4ozcFjufnb+HuHmfqZdq
YLW7UX0rMAOmuGkl8M5kkqQ7BsqyFlkLPn0W7rh9robfxiX/nx+UvU5UjIBup9a0m/HlfI3yjygn
OuhLOW+lxGuf+GyIAvIfSpROKkUL79vue0iCKp0Lw3vcp70FFSPeVGrnDT2ggMkruduU1W/nVAN7
FcUNQBr0C/3blyCjSihxl6rglrct1gIaTe2OV5lQGQbFTgLWtkX6DCfw0U8/rrW43is6njyqfWUv
gBqAIj+Qr/Ls5ViZY80rHTL8DKTw4j8gfcJ3EvsOOKCoxgPo7y38OukQqYou6vI46sdhWFQHKw1b
/zdG82d9YFsCkMm6zf1Q/OkwAnz+zqj7GTL1jgvtR7fvkgaGAdNrBJOIhhY2Tfeq3wpgIUg7ri1C
CIqZnLSNEtoWQtJs5SshARfkWTTCMYAlifA7ffdLKTW7gl67UUyZlr1ZECxzSk+Kh1tMjsbq3S41
4zaH+X77ODTde351myqNNwTTJHgGnQXrBEfDBnvlOVyHG/+babmOF/OK+bpECnvunbRON5HngsOs
WHLz5hHtFd+1DITfxoSrp+9tOTtxvf+PdyK+A1kySh0x+j87sedIBwkO7Tv9bgKzS8PHMB4UM4Zj
D8T266tc1cGa2tLBAdoUHZzBms1UoWvR0VS9sjPyeeSnqF2ueGY4Os3EXAXB2Pgw46UHGHPEQPLR
WBiSwxbO3fpZC889b7CZMofhvhnh6JAjdDtaDxzLgUorKLEv3XnBN8NVw/Q+ckfFm70JwjmXV+jJ
ZXn0DMS6Kl5J7ilWGqes9AP/fsVuXl/4o+SRGxxauX9z6IJjNG+j4Vqggq0XK8TFIqIbySqhlMb4
BYBwz4CtXoWs/M70qpY/zYO5VdigqoFG7qu2AJKhL+TbVsOZkojXv2GqAwNiDlZOBsdcPjMoYKwk
xpjdO9gWXdxtjWHVp1kjK7D2h03hn2pRZZR6nZbLNgXvG1f9Tbq83hEYU9g/a4jDd7rdx33mWRvY
vx8AMGTqk7rcJa8VCfkWX6sGmoeA8go+XPrmoFvOIsRLYru8XLv9kD6+koj8jamXiHuTDngfVcaI
4oiETTwEJJDyX0Gu5fMjf4mZWZpohmUp8NPFHYMZqHdont4l3yqHY3m1Nb3ObgnyOKpOpBIUcKo1
co6uQ4KhtdK1rp4R4C1Q8XCACPBfZdO/I9CHy/ijy9ushwsHXZZhQAYx2PM7X+OrwLrY3BPLMlJH
97M2WJ17lmzHygavq9uYRX++HEeXiOL8uHl3QPgz8w3xTVhQy5tQjHIKaNszihImcYAbo+tHJEBk
fTIauWPXQxNy30dGrk3BrHCie8LbLsxjwTXhUN17HJS7+DnA9qEQnxOhm+29n9raiPdYwsGecnGO
WrmhwIR3RC5CTSf88GtzGaKS0qCETT4slSj4NbNMIUwv5As0PyDQ2Mpgrr0dKrm9ipIziNpjiiiY
ovmD5UJOo62fqxgR70v2y/b1SJPmjiWdgk+J/fLUN3wQnx71TL6ZShrEXozI/RHigDZbV+dvpC7D
hL3eaDyqzoc1/++xY9DuoakTX6PrTytQBFjG/K1/PWJyrMBU9s5nbkwDom/VsAPE+IdtPLcBe3sR
lmuxGDpUcJcKvLR08goF+reDUpSVxqPmc1h0dWR+SnVGVPZRsqUhyCJMRErvYIMnb4DbqlpA2zYN
CEiR6qCq7/PikAIqTt5GQ4mdv1bvAOxVTBDvpTYJJRRpjAqjkW2810fLAPl5vfPgEpQRIfpJXUsW
rjpGwdkgIXSQHNC5442raGO9hulIPbAVFOL7SYhGhAIsjjqHD8pcAnI4qTA7QVnd7Ccs3LPRbHhq
4PjkFc4o8Hfv34HrrFk7Xwc8ZN4fvKG27aFq14XfMumt8jY02zyBf6Q0MdNkk9oCkrrpeKHbdIRd
M3ck3xBo0ga2YdHNl+4zIovBFFSB9i8U7vvKkExiKEHUu2eBkAt/72vY4tY2LF2QqhIbABTIk8rS
uakZJNXrjyhMIhAD6EQyLo2AYZgJSeTp5qI5T6nbQfPkmhMr3FlNIHHjtoeOYhy5NgfPDFZuC6fn
YekSQM2TjE0aj1b/tykVj+3f+v84QVD9wzu0GCcUQH92ZeZxprxdsODofAcE7d0t9obR4ejgoqNW
z6a0XuKz5nTtG46eLmzQeItH6WOtRG3z61AK0aa2F8hQYjUo1Jdye3du2A9qO+9mlrG02VSzWmtP
JHeM17OwZZWWmyJ185JW99LHGgQf5I5nGAyB0t26Zx+sjkzh69tZ+Tn9CHirdoGO3webdqj9dBz5
8TeIR6ujF6CEn1Hy9jdFZdoAwyvUzL6Zyyw1l0n7j+SZuatgXo1O43n8teFwY+TGhR+DhAdIOoAg
v7W0WxtUodNpkCRINIJTgcKEg7aeakLMb/SKGLGWZhfr/0SOO/SNK11BHjlUxFa4Q4eIe0xYCFok
ojVCe2zjWXHGRlIIc5yBH4wVbPptqRiComiBBjoc7kQKLrSIpWifcG3edjJzia+Hv16u0lmZ+Dr4
xuaRse2ZvyNndo1uBuuewHjcncmkdpkyFr6GdWUxi1wLBtq3bV/1rHKpsc1mAU5+YYuH0k1ZX674
5Ap6jfdfnBIyIzIAT1qXbmY7+3PHP8XcUW1xEC317mMovJOPAKbGfEz7XgSblumbHiKIGxfjYAQ8
MFnFLVnUstiLzLrp6zPVZVjz2RkoS66639pmHPdNnHYAUqi2eN3UScmGOMFbYUpUMyRqDto2FRnE
+wsbYcUZpHYAMe1hQ7UVD+iGw97w7GT7wi7Sh5J7+NaWWSMhEdlPeWqMhGVUF7NHNUZOI0MB8lBt
DzYe1i/57KKmGwaywHP6DzsmYXG7k4MOIXnPbKReIqE5AyCUbsD1qpDr42QHN64i7Na/yGNPlw7G
CcU/W9rZMinxZ0nkDfEW2e6CmgALIGUG7d4DpqAecNGHC8cwWSmyPfpzHDGfQGkN8uHbH8xzYooE
YH+vnURcYmZZczlOmObqzmnjHEr/CTb3nW5+nyhgvzmf5vD5JkFs1lJYYshI2vhYZveipzbOh07i
IYs39C/0vPT/mXpoZDe7Xe5+v/a2UHPYee9WDtM4mikwUEUD1qUoIXEmauEt2d1e97zBtCFitwNw
6TuaTW//xS2NPwq8xpSm5yD6t/udp89+dLBpz7VpdY9V81AVMk45M5rrijYdoSlRb+L9ZnjBjKOu
X8Eh3TtV2+4jRs2IWkYUj4uE4FqyiWp+k7ZFZPhAfga4p9RYZ7fxZZuSiBn3OiIYMewcKw1s9JfJ
fUQSGRWj5Q1hBWjRBb7QqIGFDdKZ8VMRcEnQkckrO/Rby0/z4Z2xdUw6/f3zlC5w4KC8us+aOk+o
VrJAN5vntrPYVgFOwfvgmFMGjw5+QXO16W8x7L59ytmnqbUSdLQO9seHBIub+wDC5v+LfLDBRtfA
gsIVpxUbcvI/qL4mgeeLCOPnnIxaom/1Rff+Br2sXOK2bwV/Md7SoIq10d8cRdZ0s9SwgoD0Gmel
cEuXf9bCU4Lp0ODFRzDT4+ygF0kJIqhs1IOSZwjRhvK33pg4eKZDv/utL+AkMjHYxTGpciAdYo/z
AyFHgqu8M1dXurD5PgUFLduYeKjDj/R/xbo1R1jJGNrc2I0eUvC7NdxqrUDPF5rvFTCxuvefHplo
A5AYonEBvERbW8jtyxnOYDFKBBNqDTi+L8lr0GDPWdNviKdXUTuNn8YKmHMgoRI8zF5BbYgutzVF
e/tmF+Ig7jV/h1OaFxBh+7iQjEH4vc036FRANyRAkD6sJlGKPSF4UgFdefr0gVo2Ehrbzaamap8a
v5xauts4VOst4n+HUGtSDznPm+fW66EggPCpS+HXVxS9cThEVZgCAgstt+r8UplhVAlobkQCieNo
hzxA1CcgBqbzKt5milXmWFt8EkrmzLNPsgyliCu5/YnWdIGHwdRFrveWh+6cv4cGKdPCD8IyTDRi
Lg7AeJxz5USQk+i8dONu7fiRlR7ZrRTcMOJmpM5bHShxiHxaFl0s7X2NBhmj2QPx6SMgA4sXGyCW
7tkH7kuzHV/ZjfZlfYKacuZ+uEbQPkbnl8XNvKje44TNAmQ2OmGcVxZXXQdTJvunWwBgFzbq8k4I
a/Tfadsyjt/tUzN5epCmIZq4xv0zKsbkp+H8Yslt6N8iDCN3sO8y6sIioBVZE++swkwehTcY5CHI
+ZSr66g5favuKm7nxcyAI9VXJfnnSLUfucEWnpCq5+5YN7sYZ6Y+8iyAPnbCKlrCJsKJkssZm/On
QFQNu1loEuxZK7iF4Gb+maJ3TjQvgF7ZAYP9/hd/H6eW9DnMjRscT3Bp+z1VswQFoQRIQ3RYnyCJ
R7IXqF//rYYWs4S5HX2YnCrN3wvlGxlUn6R4snio9xe7USGIvsLq9LBhbaQwWURzm9UD5OH/IyQ1
ihGOiNgUq1WBmAeAvbehKzgPtKUamB/CtXLgxPSlsKE99UnA9rh+ygDZFCdkKxJzqe27I3nQRUga
/FRPpIB8QmV0YqsFDAZsK7VqgJ3ZmuTmaXOgpWonjEWgzYhn/MGUass+zI9jsIMlRg28k003DzZc
temBznbG/05+ImQcqCxtKFGnERZbr6wgGyhRDLfskcMWVoRI3dMcCQ2cNNgrqPDwGC6X6YxHrPHm
AqCJPCeNMYWvg3MNp9biRjFtd8aeBFEecgTpst8Fz5/AdjcxADuW4/Al2uyejfrfQl/egoSUIf+E
GrafAoZfl1/kTBXPR9zFxURFKWn3WUViElugvcrSvp3fXobvu+wg6sKHEg0i2Zy8jZ9fC1Qs9D+U
lcUWz4k24jE/vW8ImACWQpCvHoLtZMP6vq9RvhtSqvInOuSBzih7XO9nyka0p+chQ4jOksMMcBzr
tGndUHi/cMoK5Pp8GTjTZ1DGZBwNxldbeqVhXbrytNYS8G1IKNS8ke9XHtP75+lQR8QTJK708568
RK2j9WXwrNAagaNujzD62wropn8m225GrdqZU66SfIWft94TTUDjT3euW6V9TIy6b9DRwt+1Gsrx
+qPQPIGly+m74vozv8iU+agfLv5M45g6PLzZUn6/Hoi7Eh+VwVdqKEoSDTjJBwNBhPtn1S7Esj2D
9nwjwtuRbgj43PGQhDrKWsgEOuk4BAYB/GQ9PAb0N8NFFMfsgwzKWwaD21iIRbEK61yRyhGC2d5H
Y1xG1ibrrBSOxwirmFERP7lcs0DBV0QO2/b+xHno7Dy6sRW5aXmwvO+pj1BKcDYBLrGKEa/dKWxd
m0cBgnU7weVG8/cL4n18B2d/1/mrW2PadKOLOBz8JaaH+8mNm+mj0XL1Pvfk713n9VFwKlId0KlO
1/kpfndffFMc7zjYYmdCqEJqZxCsr45pgaA5E55QteaU0EAUfpWbG4+vq17+662h5u0eQSCQooiB
mOh3Q35V48VTakg5cWaR6621CUCEXjtx67ZpvLgZpNyeajGNY6ORretZ2uSCKMnwhbkQsr5tJ/jE
fNe79zKWj2Y91ygIrt8/cTva1MchXxRY0lHZlK5DoNMMhWL0hpvdgg3dAOPInXIJOoW5C7rA5gVQ
63ibUhqhiexLiGbNTs3bAntuWPfwfx7zJdQKbQmR2ZcgpwzVnJBExH4/RCbnUDwp9YZevIZKvXg5
hzhpeDc4J6b/ZDQ7jNHaALj5yAOz6qTpjc/vopnl0/fitZRSxyNYZWq9wu3oDOarjJzjLMrI2PtD
iaPxUVptJZla2qxaur2G04gLWh1iW6kBm6P5tDtlFd28dnfhPxlZopZf+wQc/mNwIyK+SpgL8Hfo
on/7ogeWUAUBdGsWzjkypeO3Mka2ahbBgD162ZDmnZ38p9QjBZZBulugk04t4hy8I9sWkWmOpBTs
bJDaJQVDNxRyRrDVSZ1DadwXsy5NMmZ6poAonDXiy3FUIIdMrZ3iKnmJGKkjW5fqBaBfjOn2YhOe
tNPlSaGyU/3/E27gXiUf98DkLYz0h7ZBjrNv4spZIzNKwehs62/62vDDa7Bx/0pjt9BXAQC1vXjg
mWDhudL5qjY6vTFZ3eSq3bt0eKid/bO8nUccpzjTu9zx2BGHprTLJg7x/fzwNYtfFWnpuRpiS6qC
9W0Up7StL2eZ0mmrmAhi1WG+cRymaphzsHDKrCLk/XgVxvA/RF2tNoenwwQ8xnYFGzI6TAuxsT8j
Dl5JuLQgVPQCOZrNPNLF4iFIrA8X4hLFsz4qwGbhcdxnEZt5rsuMmgpusfS5Bzee/SdJ/aSS31k1
Y9Fua+AA+wtED3DcuFUE0NRTGT4jS1g17EA9sNxosZEvBukjQFCgY/J4mgAebEnT7HuNh74X1LoH
63CPrB648G3uMOiDeWE4bs1oIiGtvZlTJU3cd2c+rN+rzC3KMmSCRmEQeT4y31gjUjqa0BKVvQva
S0EG655Xu2Jo3YbbymN+nze+uhysL/94/c9yPeCWqgaa7+lOzsdI3o4wjPkTT+zAT8ishdlZDf1t
IKHHa0i0KhOto6VFWXjzWaR3Ogcm5BKjvxVDzlkjoUrKC92bPadQCHsii8+PwzUMSCYZdqStNwo7
mEf2M0ZD26ScpuhjtkliD+Jq4t7h5T/LhZMytMww5SoFyuEgmvv8bpYMBt0PuIlzHpZGHnsf753q
Ch+d6s+hn1I6f9U5cKwU3rkgzcH8uljtfC2HsrkqJoDBFBIjI9CE+PXo9GDofqYHrBtdRK0yl7T0
c4hC6BR1TfrcsmIt7EGc0LRCSE5SPSXj3punTuLQvuWeaScpiq4q6/1SQLbJ7k18XyC6UdZIS+w1
V7E2t05fqtLVwQQZQ8cW9TKOKOaZFD9YAMj8rCh9JgQM0gpFV99UYT2OcJnBaBFIg6TsEsn4O7bu
HFiUSGL2gZEPfXFCGGK82BipbZ+n4MwG7JAaZhq8HXo46FZh6RGGDgahJxvF68+uSIY6E4kNROCj
Z2YZMSH2HCP9XPNwDHsiupcj9UPaxCevPo4rGj3ZXr1gCylt8TPxzW6DwiU2CuQoiQ41YjG+USHx
U+nFDybvJ8VyJTIMzPTlhdZSbUOrWMq4cdB91e+Egcxfal0eCHBkwIIItKAE1pEi2NeXO/pq9219
JipTadOH3ZqkKOglWk/w0jNbCmxg97wkeJl2nvx2d1jvDY3UkvTiEGnhwPfTfHaNSStK3So1jxsq
fky08VxfVcE4rnWBqGmx9yAg1Em7Ya4z7n6DKHUDz0Y335BP9L251mTT1G7r+HB0/e2x2n9dr1+/
SSD/ZzbDCfNipk9/iNu18H3CjggyTSnth3lzglEckXVxN3yEugAfyehLHho4vQpUwRxD9sQDVd2k
zNB97izprglfgJg/BDfmbik8KRyQl+TgcN04CyaadFJ8LaAHppc85Vm3qSiXI1/1bPh+5vhGufAt
M67H1T70aTS1QcVmHOwA+1g4wzWXGmWC5UMMcgEZyfAXULiehMa11hVsePX6IVhdUEAr158VJxnc
DAX6vRDZCdvw8I+dAAhWHCS+8QOTQpfhSI+kzZUm95o3+JbfFb72+zy+1SB1+cY3GYNXFvRWEdTT
di6ej4zCJfdpc+eM/tba/pQ8y83AR0MGClwmkZLcs8ueFNhIvHae3e7HTFIvX4lSy7GHlb2G+GQw
lxmcc3HZS3QbvJWvwm4GVH/Cf8rnKHSqEi7hVCYxIjDpv8Mi7zwxNYZqQG3SoJpQQ9/H7NB+D7Y1
DM3aETa4AtNbC0fHs3JgX5e5Z6zBM6DzO5XUeY5+m7i3oSN+QfZXA5+I9e9mzaC14XNsLKhPNhUg
kvty+thNuyRxrpWKnBvDnoeqU+sjL3f492h3DcqbrYZfG2FuaWGGVcCtcLT0YwK/Sj7RPzbxLOFe
uRznA8FztyKG4NTg0ezhGeVqHVs03gfoeGUhD+MhzwtFvEUBaguVFkc/1LdkB6Noq0Av2vVm3CAQ
WqwuNWzllIqbmWTdeJ12n94LIaIT91bSRL6RLbmBCtPB3MSpAFJpxkkgMRTLeffEUFk7cGbHmktv
GMvowz5n62382I2dhljucsZ0sX6KHoTnD2OcLL3g0IAHticNLQqSSr3XeDQA1gQSOfhYQWTcxI12
5dJ7Giu3NginGZ5vUGbE2P4ziXoK9tR4PNRviuoEFVQpfHeAozD0DQ9T2MYpphFKhlZZkAGKaDPu
dUqufq5PYO3UTSBQwOEnyr0yCVR79Ba8ajeaLGiTV/p2bpt5CMiGZ1z10FFUlvkRe/KOHN6kd6Fo
WKFx4KbrIHV67bDC3CNyK1uXGfyTHLQyCMqy1NPwp3ppHGelD9orf0A6eVJaaTBaGZxPY2gkIJJc
xnC3X9mAsYjdGTVeTfiNg0fHKR8MEtex7gbPf+sdDn0Uc1Q1nGzADlov8yv+m42dmOYSQ/1tG9GD
Uzbxs/JY+iEhnMxRtKtYmp6a+WqtO17EGWdHEdmLh5bfQAW3e0K5C0x8LzwbicRN2Pl4cbZGTl4T
ai1bN+Z4A5L2ckTnF9gEYN5j7S67CoRmvvCssOMqwvBi9f/XhaC3P0KsmIjoOuUqm+WZJo3RgYmB
7zYwTyUyuooQ9dJ4yhjJ7cBfwMQRfccLf+C/ULjPX5V8obFtRXxfGDKr2w4MU/SREdcaElKFflMY
aW2vaQCNdvDMuwdYFb7zRUmHLk6OznN45YKNQTpd+hNfy/wePNjtzG448Y4SHKSRx9MpfRH2kPdm
il4BoCIqjrC4HhmvuNfzoBJxzsHgYxthGP7TWeRUr1VyegAi2zCnPJPCMQp78SpJcSdJZIraC0OY
V38duo8rxCAdPdmlSkpXb4cnWj8XA8i/3vLQtDFU9aKNNahU5TSj8Ph0pzSe34ZePxMbrAMCrYQ+
vZ74pmu3jI7V+CPFcAMDo2Em+kFy0jkDgh+Bc/CTbvvvciU1jXBTaMldjdDxHZIB+Q62ZACjzJnr
kfuGOQyMpoiwb/T3/qO5eLVCiVIz+L8gvSEghTD09GFwuocu9BpIJdRbLZ9sNLF3OLB/NzB4VmnW
VZwsHtEdNmINK7eIJ8YUT3F7O5Etrpdnx6NkJG302sROdM4YoB5ngemJHbEAv7BV67OEBDAJvNVo
EE0+v5U5OD8Y4abo+xScfE/Nzd86Kr76L8j6HBZboMPNJqSHFgq9BMIMgaoZu38aCSU6WsYwJyPg
1uCRbF0oAXaVX+duxUSCdvDx/HNcmgxONGQCod1688MZZT8pGEzUZ0UaA2/xs0499pAFeUwdI3Vq
qDrb+7cvkMdEDgskDd7xGUtIIsJ16NsltFVI3ht1GQgEr0KPRs7K387nqRa2nWxRd5GMDOp6CmuY
Jpgco5Ttu0GeCGtRAV52UcIgtuPnfy2j43eHTse7OvUCXOLhljJXtnLvk1ixZw4ZCSR3P0gxDQ4G
r+8xjUF8Kvk8un9nZqwLUWJMi0NjdiLFt4kgFUBXAN1xg1nApZNyvHnO9DDpVm60Uz/9bb7f3Pgq
JRrCF1dq/Kk6lxhO1YwdlsdKbZc8m2SmCr5b/M2X+lKKPhKiB9gy4x9pLcZoJDP9vddH6kTq/e3G
iZIeKqhK6VJHJlBFco6RYRrcqqC97QsZ38Gq8AfNIVtg24aedCL5v9BRKbdfj0m3yyt570+b4b5V
1zNbqjk33Vjub2p9GRkgstiRUqYDvNaVUi+MrCVpsjTo3nAv75xP202FIA+iMISErvzgTrQgQ4bP
kEvXK58UEf5aW2CXq4nkJ51mGSrJlwhM00pvPKd7Z8c+au/W/IgvjfZUAnS765lAtZRM3L/JlFuw
rDT77Dq+nNQF+vVpYXBIevjWDPap847Et/DKPAVadt+mqgNUBbGyIOwYQqjGwpDDCAbE9quGNTC/
KGSj3l4vN36hEPreeR0iwfrELDmBJioAE3b9mM0eUi39N2YB1kqb6DZrV34yMYGV9VgyD7qANWG3
FgMRA+M4gIgLJZKLC+X9gpDPxqOU8YxxXkWrUV0YjEfyxYm8KL6UnQXpMpBK8knHTgHFX22uYFQ/
pFfYAqjSPM3zWFdgodVm0FM2iGx4S8ys3TFhuJpPTQVa7tpAvn5ep0ygyum8b+c0tuEvfpXqHzDj
93qrzYuxbZmUEeVDq5dA/T46MuLvT18WqSmxgBRngBKOwphqTK2dC5XyUHUjzOR2u/QDbKP6+9bB
QYJllrML+TURj5nl2FF4r6+c4+bS7DvOcUQrK/VHQNstfpN0AcP3XHpCtrX/x83BafI6Rlfjo4LH
Vd6+VtbJU1muGa+Bfa25HPg8rErH7nKMGFh8W4G/gqHPRRf0fwk5O+TNryUIVqXcVUW8fDGNkJ1R
c4AVsr9z4xuzJ9pEuf9urEGj68x0da68cXlkyMRu3noiJD+GaV0g22Yc9L7FNrBN3HJVNdrmSYpF
RiWCrMFkmliT5CmzoW73XCGUlaRAoKxWXNBZrzx5Y5MegxLDJGQzMozoz/LICGm8OQMg0Gc1Fqu2
iD/BWVgg/kmm5zWsOc5x0kwBYnxquVq0qKi/ne0cyL8ThbEoFxiBCenwmgGZl1aEdrK1p5ZoE0RX
lUHZ7YMy6wUIR3yPWRC3R5oU1EnU0yiDZn0cYnUmAZPq/M8lNphqL9kGYFfBag8+MD3BMeMDZ65x
OY5+6eV827vtCVq5Cir/YSY0R2C6fnEWz7rbVITct/xhyY0I9apkRazAZQPFbZ/0gixcJJd8B9t7
olb6R6Q+n2tcUk6VeSKhywbkRuG2fNSbxaWXn6MPj1RLxXrO19szribtHFdTm/xV9vdk+08SK+Py
JV3N1mGmULWEz0W9B7jKu/RPjxTsbNt799clBNLK/UCLTLLtzeg1bl96C1J5mWKTFA5QXHI4KnY4
CLkpnKrYtJQQlyk7oLrQ84jvmIPY8hV7J8mo8roxFi3wsIYJe+7BzR9l4YJ/IK/YPEYKVhPS/ipc
/YiPTVyC+DQvsukingL82eFnNv7NyRKToy1+e1+A2C2PZNsR2MjXLJi1l3AQjTNHoAGVEywlMtZp
mc/++PLnIH5wNHb+yxL+UYv8rsMTwz0F68Nduzp0SyuW0PQHAweB+ld4x8REuzPeXXlDAlbalxSb
BOGOUkvCtVYtGxmNQtmhm9LGR4qN+77HJKZ3D6QqGNCvEp+OQ91qSipnP7PtUWiNW988GApPg/3g
QtV1ql7msR++Y5D3JY/q7GdPt/h88DgzbJjOPOngxUr3F10CttGEVS90w7Vp0aVzu9BEBNB6lyFK
a+F3z7PxSmPZySZ8cFAsErLt67peTtFqa71mIh+4Fk6d5XiSNjpNz3z/1CDJcVCzu+a3QoC6rg0u
33Pf0qhY+9a3jZxGzZq8OcxIzZK0rDRlF9yF12AUMQoqwPfvspRC7kz5ZEJNm0kJaLehep547oKg
VG6yzj9rst6BcOBa0Ws7jECI1qkIfRbqcpZsLs/n1Kc8Ah2I8uPrYdd1IXyX86bZ73Nll37s9Y7v
PIwoEfP0OHYm+6pFDGL/wdAmoPpKdBXbgHY3rz+taWPj3pHIn98k3U/0A1pdDNMqFuC3T2chrAix
AgReTeNh00/D9a0Z2IeCC07celQPNbk5S9kQyxJ1uXo71uO6Qo89ZcD82KwX2cujYV9/FoFjd4+Y
zj4n6cp2/lLxxOEwPXpMr1DaA/iU9f+8fh2OouA9us5R81v6R3QwwAM8kicBViH8TSn8D+arrkLn
sfCarsMNp8SfBTc5kYTzvcRDIFyo4AH8w2faDSzSu3+0BWKOiz8wW1mEnZ5Pacj/Okjzyb1MDK+l
r5JSqCKOqsjqHH43NnIuoqAgpTOHgXICFJ7SeGOI0Z4JJM3bvQ05bh/MO7qexQnarzKApW2uUs6y
LSwm8H7aci7xZO7IvOXzEm1Jo5tKf9t7Rhg0V+qj+wyVsJylHrC/yIxvS0d0zvDmDNijNQNjkBT9
baOkjQV4KlBZT85EPB3BkZ/RYZg/TyVqLhnsv+8Bpu3yAp/0Ywf2ziCjIJvbKjmwccha6yfLMpha
IO7x3a2G5nnaqIY2LQvP2+sZVRaW0sOdF1IPsMTYVHE36HagBBffSs8xFft/NIVxaEqXM1o/lAC7
hL3biVGyj0UFbNL06lGppE3wCmW6XEshFT8R6nc7K98FzOI2dYrmAvf/aJKsQn1zBreLyagXx9OI
zzX3QvwKSGzFwCq3RXfvNjBi2aMBFt405w1if/k5Op+JJwgKpOknWokAtCTzm+tj+S1sTnXAwymz
Llwqds1PARTxd1Ilv78LLgzqI+bdwumVFzoJtW4X3F3ehpdazvlbyu+qRIuy206/sY+CWf66JPU2
5F4yP+0IKX4aAKyJiquGiezKEWto/WAnq/CpLjbN921AuvlgVZIIX6b3kYcaO7bQnuDIOx1Vb/pi
jkbUV19Xyje7zDQTxR41HET3geDfbjOp0RQ+pGKM/i5SfF6SnTIW6UdXtGJpf48dmzHOenVrYcaZ
lwTo/29xPjGzNNXBNpaTE5oHSOCcpls0uIBgOlEbQlmKwfTC6voNu0fyAfKMXhn9jt4S/+pZ5Sq5
CfCn4qk4EUvrCpEgR4iZW+lD/sRM/BVOjTE/Ej0wAJgvNjuTUzl5gnLuhRSzSjS/niQWeH07ofQ9
bky3BxYWQL/E/nyiHc0fF+9lJ98LnPuDnqJkLZ4JyKUr08pQtXxshepVaoUpzZFPpyMO1z8cRyZM
HATTe9rug1FH8/jj0/jlujKpRlditM3VsYP3HDd8uc8HWZqZfF02TlRQN+N9c0GRSXAjQyv6YYm+
ob2KBc1bX6R+OO0rSB0yK71WqBmRLj4u0j8VmdaHUNX/rp+Z0zOGtN7SiNKa/JYpfNlihG2VR1MK
pJl+WRTU7l8tcADBOmTHautKy0KNW7LtHH7FgwlkK4mtL6VLTpKk6g7beBRkYBCym8c5HiNaRLyg
EbcPrIFuXPP4V8PrXpQu27KhAZXW+4MY5iQ1FEIqs5LhVZHos1ohNVfeFnHbpDGMtycaq1y7iJ2Q
heg2XZh/fBkQq5UAMDzERd5kflkwnF723MMKp1PrtKqdB5ZjrPXTLToklpd8U5uTh0qvuxUCum/e
ieqzxYDCxhq4IS2SmGuRGgURTN6GLuVuGAaOlULc0B6mt61NUcTz7RgYu8r4Nw0qpmrOSbEwXtLe
ftVS4GwuB52FQ72ahjw2HYUkcp6lRiqsxx8qTehFOIYfLTKFNLUGuawz0E2LIJqKKh2LFTvFpJDq
kJ4V/reovXmvnTtPBj7OYcX8dmx1jHxWByAK8VA9UOtsqlTVcyyiPcqMf2O7AkgKXEhETOmC69/R
dBL7QSGh40SqK4/nDrOdTLBDM0YinLFuNZLI1zxJ5xkG3imRSUx3NBIYZX/vRG1G2JE64S4yuvA8
7MX0O4SEUXwa1iHE6Dzd5F8elz+BbXcv1oOc+8F20O7dkAjp1SOE4Cg3K6tPMSssvOGUB/9SCaT4
zMI/MZamfYbBCChLYlhVkENak71iNcVTlZRegCKD9YegrR3cZygVRLFSs3AZjiRDLe7VviV75+Tc
Xkz9iZbmSCpE+OSK8hstVuWKIwhBlxPcLroWhaqpiHjSlbroMMsiASKJOCVYc+XXvwSruUPenfyb
Rr7TxIS4PBk+s0GQ0h/08B3wffjUFUb4SZt37HURODABJ1ZXVJvVCW7w7+bPYt6rJ1KjBCIkIjdj
tsBVPCLwwdwxFhgPq1CCel4g3HetybsaN+KeC0m/lz4DRKZ2mFIlf+0Ftm0XgyeQsSPTUGd8Xuvo
btu/r7/GojaemX5HWiS2H86PqC9vZ9pKwU/mFTti30PqRQPF9iYtUuTIi4APMsCYtDPtSrde1MId
L4ZDcV40INwIBm5UlHz1UDRivz4GRWN5QBWfoBmDwZaA2dpxcpiOBj+0rKRbuDhBAUsoxME5TpRC
Uoq39sBXjJRrg4sTfQy6wC0fvkG09Zlin33qcVQm3SaDXp8Q73LAXUV2N7JKBsa1RGiicF1xNCHf
QtDmrcety76PF0TxeF9OmoSsl6/ukanGOd+1OsNCUW78dNdeOOxFL2T9gvB8W2XXSyvYmloXxH7A
/zAHqqw+2MZ126InbIlV+u+zuzrhdgg8h4toNuQXnrz236ikeRpS8eSF+Bdb5TKjb+am7jiHRrdq
GsglIoATb93XZHDifv4ELsfTavuGpj++OwD3LbRZTd/WFlZzV8jBelOiVnRZGbvQ34ItEjVyIo0n
TsG/pDSkdnWYs41UUIogEmTCOGzp628j9YuoERxbFray3UmKD+ejoO5yQLvtMxCMHMvsoBxBI3VO
xEv906DTAL5QCdE8AkllSjX6qWMLlNtGYU4LX4cBmk5xsLifWAhXTAMV5kggrI9OSmQUimLywAiE
pE+TDVtqwUd9vSSZgxy5E31u9P90wiQZUHnDZQA9jm5PqhPoU8wnLgM5JWVuPTdGXfd5gZDA5yDG
wwgOqIlqT7tg8mlOyZWJJIYDawjdX2i0ZcoVSPRMdUi2vb4pMEHNhrPOtMHRzIAAXRTc2yMyb7k5
rD3e6lB+NPpgr6RWVQ61ifBpsb/A14a/JIkinNeYgfxzlBXTc4P2IzRhU7obwacBKoNK/9oOXZQQ
7yBnM5fNt/LGfv7ig0ad/EDj4ZIZPQZMHHqjrWUtB5F/hUHHwsfmK6y/menGFH9FsFRkMls3w9K9
elJpZUoZawKhWf7pt2U/RnLBPNLY1TCdH154iVx6QYSbKTLoG4ytOTHGSOhyYY/UnrlLKPEimpNC
jodW1xwh+V59qvS2EUU83dj4+q678+yIN3/jF44td6SwKoVGQkiIHB4tdzChlTBpSJ6bADbpTewJ
Ha4gnu82zQRKuGEoREHS9FyqtgyMMrJ6j2GXIAX8A/HT9Q+VxLVxQY32DhXJSLFxEy8WxSxPv9az
FsJQ6vtX0Te3N9slf5efhPRe1aH7GJDn07LVA/S1ALSblxMAPw031C4otizBHXcTx0wgTYjszsu0
7vxL3JDX7ahKF6GYsTDFRuvM6xgPloh6t58jaekddDxZc0HnNX5u7stvUlI/zIoSajbWPl9Qrlsb
k5Y64vi+EaPlKx2Nb4tyvWRa+kTuW9BXzaWjaUq7M1TU3OrHUfTxymV2t4BkgeVhqN94zgQivrSf
k09K51fN5U6hLBtfT/OpdtafRbpYfB7BUgcAywhuZisXhhpPI+pwOx3b7EPoqtd6MtqXRuHhtfGy
MKUcHRuUCOmkUTOvetZJYxNjfhsMusSZJZEOjM+yPhPkxqizu6mg9jwOfQFE1IKIxUYWSsVGQmk6
BeOLPR4dUOyb2SEDEkSQXk060J4JY+xeTyIghPw/myS3cXJbRcnW01HMu8A0ZFnVXxViHYrU2vTD
bHj7Egzw0EEGr9qEBOkvuZO+QWsAHRraHg9tzs90mI9LgS0gcR4yYJFVBLQhpLnWsk7x3ngA0BpH
55HWKnPsuFkncCjqKDkkkmKwLc8MUqgrVSYWgdLMTzg62v6aNmRGD7IGzTiEGujkIP5aDWgAHueZ
AKrq1d1XJLDCqv95PCbp/EAnH+b5A5goGLXf2ZU7lLO3S/qED1b/vGR24La61YepPnaoenutR2zE
vto1EaR3qKYopUqSS8fg/fbObE4TRmT2nYads6I67yYkFNXj3c29lzMN0rrWZXR1jFLmjFd10l4x
gmw79pOGFqNDU1YviZ5QPPqdAc5ZTw2KjjmSYaf9ij6JgMx0TsydakzmAITZ3nNflOIMO7l8DngD
/eV4iKJ2OHhMsxaZHwl00RvWGcwKJVR2C0gAFD5Pm5BbT+jwlcZzb0z5P/wu3S3WbRjaUQ6maUlj
0n4h2rGUjsdpFyB9afnnHBHIDa2nwwsx415jJTTayXCezyCyjgr+dftDqOGrhNGjmRxRIGOxwbc3
KrGe+1xFp2U2tXvD9L8ZvFT28Lt0w7P9NNJ6W7ddO//2EbQEW/+nRdCRXtgLEoC5OgOcAF+F+gSB
eA8AfsL/45zH2TjqPu3hL4weGA1Ubso2PJrYLPBw/wi9rcWCKtl8RsPKkYcTR4S46haHKAp4TLCJ
gv5DB69hcNZ7QqbHSVnYyRkl7v3Hnr1vQeccOLTqp6sDLbgZJFe0Qa2HDZsWe3CZkuh1eaZEWZdV
yB/EFh7WnsOSRRLUEsIRy8RVSKLhm28Ta+AF5oiRdvcX8rDt/f253zGav3QbzwialJllvISat6Zf
2IIzneZibC1ZHBzHXQvUXTrL/lWNG8v7vsNcSyHXJB7qnRdPkkOjS+wwJIdS27DgF+x+p8L/kpDo
C12cOzGUEp7AjxDrWe+k4flOLbp3bqkIbLigk+Icf/BIKwmgpe/WjcMvWGEMiYIO+Dk8Hlv2KxZ9
4rB1jKrDbrgfB5OzUIrq9hXfWRs7+qf5GbatqSMgyF49hLo5Xpthn1gs1saGkqfU0I4Mz0lFJY7O
D1EaeZQjSVh+Ca3jT9otQ7w4cHDlZnHOsO7+ppbpVm1kWeC5J45fxsifN7LYlhn1IK2Lrx3Rwd90
9ioLQsae4lHuLwHaX/rTMOwy1jL52+AsFGwW37oVsQKUOweP9mRbfPnCh/wIziCSmRHsjuLfYkz/
32h30eoHmq2nT+nzc9taKPJk4tcfgQzZrNIi0m1uPjiFyuRRDPEMZoGp1CIZKtWvyLOA7vvo3vwg
91Fg1sDp59rq+tDW0bSe1rfzxIsqke8JAoo/6WQdhKDI1r2JXPsX+M78iDMTtZGBZ1OTO66rjc1o
z4UjBqnYeVaaCmOlKlpIEJelyhqb8GMsHWdkdX1LSoiDxqqd6S56VLTx/dmnZRcNd77DY8wpnJMn
ojvuafWWrYT9qYHffS5S2sX1gm2OA7zl3jpJAPVA80QqMDy2rPJKiyGYLgDO5YxHkl58alpyVonW
Ge3bz+vtzkzXqbEaG6rBhT81DszTMmpbR5gze3z+sZ2/6Dwk8j5/Woj/uSLDHVGGjwiA6+kFShV2
27b+1zeH9YmzHJDavlae5UrD0dWmTA13DVqkjP9DJBa/RgLSKzq50Esqf5HEfMrIeIfyxEaPKOcW
Gca2zZiYNpwek1aD74rgXM7xJ5Z9yfnWkCT8F33a//bFRpa/PakuneAqYm7pFAtwPnw9vgO+HmxZ
I89h5r/81oZsVYEeQCLFR1CndmEmV2sJtIO0FkYxcWLmaGmI4QtfaSETd/qSCVMMAIWCWKJCoYuu
xLZQW8czSVuZ4NBBMNmbXw9Qdt7526Bx4XX3P2krcU4eS2l3rT4fC4YVW2tYFAaH/cJmJMZGjnV5
mAdcBqw1703AcAn4KgOG+ScGYzyKdwmCAB5Ep9uJOKFIY65lbb6vQGpeaeRZwus/Lf/6JP1pnlEy
czvl/fACYfbSovRnpYFRQP1i7t7/2unr2N2Uf3oFrQmPXkzVIHJqyVqwVAuPmqGU5xiLV6b/WO8o
ZuATgXfEqPMYdgTDVc/lpABs7pIgvcJFPH7fnaXvKVlihVQpb4XIB/cLT8uS978EST46jBAHtQyW
9N9z7taCyUJMeuK0RBSiVHSm0ZsP1EsDw6Wnab3N5TrOQc/LO7OGwL3hsByKYMnIxou5ls31eH9Z
1NNYdgVd3lnbJXO539icU/E64HD7iN31Hcy9PfWBdISrqoyOGWyN5X9+qH5dXq2+KuP9DeeGFLur
piMRJD9k86fCgHcTMvrF3WsRzRZPsas/oZyfIQhgAMg73bHEINxgAp5sm2ngUGGux3suGxFQSdmH
nsPLa3TS/1Ev3XM4AGjbTrtiNPVQMzdxScVoCuhIx7Jce3aEiOWq1gRwTz5Vsh8R3cf/2zvywZFr
HoYnzI7efkUgbH0Nnmb0PasGh4RJuqlzxLdWfakDjApJoNLH/C7zYXUl1GhKLC3aTqBCIIeg1iao
EJWJX2JrpdoJzVftDaf5CBgU8lEvdv0Vc40/vzI+leFPeI0k8VJ6hsRYE5HftBsAvXBBPNtYGLg8
+Ci1eQiBP9gUgi8mVAxBNBHk7cldbh/sbCtRV5C8gnx3r8KWyZauk+waTxlf0lZn+6N6og3g1/BW
qtn8ctsLfndGuciARvsQfJmij5yckhQBOKtGhVBQ4kcn6oBzjQnmeNff3cuuefDrJmmHtWbEXZgW
l5aJmZ1LRC6c/xX5w0FOuYDYQWFB4zmp/wnpyXa2Kg/QRTwEyBQ3GrSZEAX2goo1+upLSFJY17BU
DMOq0CqfsXc5588UzAYvQRf3+Kyy/NY3+8rkETASHhMOjP2dkR9LVLn9NdybbSuATqvUDwLKQu4N
z4++kyeO3r3KyKTyhOHMdEw5phmV2+v5/7dFbUdqulfc+2JyeNXx9pK1UvguTiovjxMGJ9MmxR/W
qTt3+ynVs52Gkb8uxYyshG36z5AwpMc006wW/KRzYLCeddM/YQSCjFiQHjdojBMRk3PZVYlvjoCC
u6cSb/R3l3M9zRr1FomL8G9yThfjqOJDDxgIGRyLZoUUotMpLbvEFuDwL8ymMptI4QYKsaKAtBOA
c6YqWlLSH57esMR+ZgdDls5eh5XuSe+OptctsDBNh+/l5okBgZGvqjy47FLxz3oVFpbcKkxgZu1i
px9vqwvvyOpK5m86w+Ob/mpqVXLgqpiafDXwm1VuZF4LThX7PW52TflgbICxa83C/QdUcf3ilMIG
CiAJmo3DEIEDZVhkaGdJM2Smw9glcXO4jx/qh34zQ8QvEC9ByCxma4XUgIm1js/vjCnSbuhnW57R
ezUNHfmfcVD4FZgGtAPUrlbrJwBcNnQT0ort+6qlSX+HL5t22S0+AF2fYEBTtNdB0IzqLNwYVPRf
mOzh0gUk/H8hIp8CIs5m+0n/dII+bQtgeThQWefoFXl/FbzXXdmaJFU+omYMZkZuBvUqlUqa2KQ2
HVUR4p00C694Hgh9Nix9gufjJwgWS6JtMoaWZVAXJ0ORWnc1bOyZCQK2Ow5lrQOdi9qR8xVqgys5
DsKxIdpw8ZUiU0kZZJ+Zmdj3WM8gTzrcJ1r9R1pKm6YBNagYhQMksVNMrtJh7eD8mwPOftn32JSC
cE/IXB9ov1qis94Zc9OdTBI0sOzrfV9Yjd+lIgbcUKSLRJyicVa3gyNOF1NYF0TRELF/b84+Xhd9
fBNBqivYHD4P4xerV2PNi5yAnIV7Eawp4luTi1UYvPAjIcUMoziJqGFdz/GNumY/6DkxW/fI1RGk
syrDJayq3nFwOSYC+xGFeSjZM3qmeb8Nl7Ym/6DC/zgA7RkzbMHenNKY76//G7fF84S9uIlFYvHF
ZCGlVLiBvuCsc8MDXbHUr5ljhRwZUPOh00kMtbdnL+MdCzzLv9I6VQJMas7AH1gWaph+m6EWJhbz
Jsbc5WQwWDUhQZGR15DNGC5BPV/cuDEziQ8dDXUfhUGNunfVSZ3b7rxzWpNgNFQ6ugkTI8xlkzCB
mL/fwvlOdO9tAHGQt1/mJae1XvjwUUK34FLbI7seQnMOM+wrKMZIp6QLF44nYyjfNkN6pSRaK4Ui
yTodxGmNcQeNk88R1/tUe0n5rVFNVRLxEvRgwdhfNxgzejSQXXJZKtJixiXlEKEKh9A40BO7K61i
lDzQGcuCmYQ0cKx8mS8CFx02ModAOi75meAorQq9Y3pxHKBHLhyZ+KvGRYMbPj0ZYCuUNT4a0DG6
hUPg2i95cSu4r22m9+saPYAjhLJDnA3tlylckOZ1BRsBHA2xh1krba5TRb5IEBp9CBIh7cTVIRwe
oPIYA89FSbATNKzzQSUDnvSghjvTmbPJktS+uBgMZrMaSXsQRL/SXBXPAsBjw2PxBNkp24qXCTZ6
oCvu77vEIkv/HCeQJ0nYvgfPSm3MAgQnRjwvOXBZylR052ohJqANalqrFbvcazXvKG1ert2N3nBo
6Nn2kNJeB6dN/f62ZRBvOP1+ygu/P61goXheZlGP10iagf7oO1iSDoyn79IEBeKMUPZdJMBOdBdY
aPZSF6Mu7D4fRMJzqlGPH8yI/L0V7EWBXiCtwq5Hgo41XxSDNQQ1TFBPfu5596EbtR2NrAsU5DrF
DsLDXX0GSO2xOhhHhlkA+ToM8S+2eDxvoUeEbkHYxGtIu2RCiL7xPWWovxtccHlwUgS7NNfVutH/
0iOOG60eo7LTvZ/PVxLgnSokKx+q5TuXx9s+E0WY8KAeWE9PexPdjW0vi+yxd56jjAzLXT8/oxKm
zdIIX1oUWK75p7nnQr32oaqzY+CdcINog3QWTw4yphNK4Uk1ovPAsDqitMahca0LhnxQa7JSg5qw
qTq3GkVY1XnWl9cDmsymLZXiGGllaJGQCfOgL4dWatoPQW5oaJwSi2yL/64Lw9CfpQ34VKkZagbZ
sU1x5dchFGbNXQFwg/rfwFxYlexP60LNtZyUVTpsxmtgZXsRs0q3HdEb4eYxL2AbgXHlXlMz9B8T
HBUnki3QqReiQ4phDwaCqx+HlSrMvL2nHyLmkZN6PEqP7EyAnfRgxcxLjYBdG/a6NioXrTA853G3
v6HMrC6yu49ee5EX57MpavFFjGwTIxr6K5Nr8T9DOoVEUM849p0GqilGzJN74xwN6hxY3KYFIEfW
6XYKGtkVC0ixSnyUTSlVEzaIRRb/16YFayrlK7dGwe6TbDqkYyDfGmphpCIqhgQ8mLr5cYjEBCFq
xrT0hNmcTia9giH90B961OSYFcvMgvvKUy+ys9BjT4Vakxq4PiQ8Yq5g/Jm9T2EJLeeCTt8p/tio
MtjVnBtH76ie9M3qzMX+1bG5vplqsYqiEEtAk0RB2Ngts8gD9wmzH5G4JLhRB7twA6mxiC6EB0I4
lKA+CpISf1IF4itb0lX/T8j8d3HAz4H9pzkf183yOGauSp3BhPLjExyMIduwMteU4s/pMSLc+m4M
dI27veegEBcyDjlTQi2KyewfjhtLQQEg+AIrTiISIzi4Xdy2EQ7epppykAx+3OV7Ax/fluXX9sVP
og7hZUTeLFy+gRTeAR6vw0l+SPgzAA3RDqxbUgJAZvwkiKFSSQOpvNH88oYuk8gLsaVot/nJfDh2
2uawIj3uDRd8krpAik4cJNcv1C9s8hOsnexvXunLsgx4uZZ70pqRxkMbxWllAT8dW4tEb2Hf1FeW
KLkp8ok/DeO4pITFbKKQkKqRqQs41CrZQTy70EWONamixw+yqPREG52KLSJC2Pk1KfxBK3M30S1a
8U5qQLsKx1zs+Az6MRHlCz5cSYH+IFY2BRqmvOkxVIUscVC7bQ6vOsTJgQ32+PoWiTmHLstw7CH8
mwtdVhrVTmbekjyeHQsSMyGpOmFHpwNlST08vsIFFH/ec8ssLAcTNtHfwK1QDkNtUsAYPS8P+Nm+
vNEfKj4ehp2Y07zKlN/HFa58GM/q4ktB36wZGwVNaz5Xb3sXM0QhkvmZmv3xOqyABpG5bpAN6YyX
xmBJPnogBkYNTrG6gSp5HYrzeFRmCqdRhOq7eTUFSWRd9ncopkpValWuRVIoNe9AXVYCzFw9dUhl
LgO+byfj3MW64aG8Gk46jar/nt3h06B0OObzN5TBG0ytsA4icnMzw+jGJN4XX2625U+eEuBGQObK
JxW2XIaU6qYY+IoOikP8f+ufHxWEdo8xBGYGdfy6XoDBMLSZ/b5ZKv8bG/4rqqJ7pJ4prFlaFcs2
MzrrNs0yiHDlwBKJGVBFvJkF0XhyEmwoTKUU/10ixu9iT+CqKtQ+DZCZb56OVjbL+pxLHk23lyFL
DGx7FqN2AoAP20q4EHcFtzOclEcshOoTjM8LLjdEUsEWEeYdYblDGv8gR77VnOKFawAYm80IDm0m
M3uSujSDfaxbHLzrXosKF/GAQqyOrDg8cuUWM4JI2MHKdDMzRBlPkdAfhwJVTR2Aq8gg8I0+bHSJ
UeE5kABuF59/IGb783oKkzdw+HPjOyDdEHeuMDV6DLr5v0KRAIlV2AEsktT1U2PBf06f88fEKnCb
JLuLQBTTZn7RaV+MIRZRLBhixjRsekM+M4oPrA9qwPaeRwSqJjE4AopLL5vk2EyvH9Zgz+AmhsIA
6xrDTUUsJyUF0NcnViIGCyTk6rOy+CmNCwcDskVna2cPVfIW0+EbBTGBT2ESXnEH1dMAiwPHQjhj
Vg6Xb9P3iaovPdF9fJlG92RhNBE7hvEG2nC4uKpE8GLsiLyMQ2Mp2g57Pe7XUhhvR4lM2DWU1Pi1
zX/PyRY92pWchNIJtvO8qITzqy1zUcU0Yk7anW8kM/96FkdyYzd6m7NQr1oqPBNFLn/FbTrNYbIL
/WSQPRtBIOfkM5/Ts+zMnYFED6jTj422mI/NiYg6tkZNKsrvXAStnUANVmpAt+XaMpHR9CcWdf06
9X8/GFgH5rrrZoWtkhn0Ak1knmBDFN0cKY2aeCxn4UsfmlVhQvonH4zLTqe17D/Zz0+hgM7UaJo6
Y7/+/uum/mjMp4I8A/PoG2DpyiTZb0GNBr8DnBKulFbHmT+x7DaXy72UYQcDFgZ8yiZeHcVwffY4
BD+60hNIdEGQb5hoA35Z74wHx25tPXJSwjL38IgqYdFtb4BxfU90SbZjPHpsIhG29ibNgSKg2m5R
NqH7xeKag2rPFmukFReWFDMQfipKaGku1EeIWdI8mSI2cpZual4dWa5xL9fEUKzZRtpSOJG3AC1m
aHdSmC6jptZZVO8GoGKC29h4I9+ho9vJkM1pji7Fhgcbsd76z/1NdhkvW3Ee9WC9qusZEzFvI9rV
te81AwHiH+tQ4Q5YiMgXoJODh88rPpqqr0p1QnYRiXdiChWKAHfapQxqWOmIsVhZZNXWpFDkyfGH
r0Y/6Og6T8R2tLBJZBrqui9xULyiFobm8BqL5mvQEnWmdMt4wprcXcF83RU2PbsAIH2WuQMJcixg
dACPFNOySweTJj+B3f4ihH6oiENdEPfYot0pNt7eMMwufdt604ed7p6hCN6ZXJG8EuGuZBN9myMG
v3mr7sSLe8shnUNytzt3ZDt8Uix4I0fjVzUmlT61VbQzc1eY4JypCszj9SDzhmPQVrv0YfFsCtLp
DUkTpIRmnLFE+VaF2iNkxvudJYd+deX+jEaOdRRfL1QAYXd93vTCkOdErA17ZxdQKgYK0w61Zh6p
RImHWqANN5jxxxBcLHflFbCW49P/jphq3h7oWCLVYoX3EJKHE+VJ9/+YsyZphhmZzbJKx+87HAys
T/5l1Y9TTYtWYSqPPbBNGDwt5Ax5u4YR55ti/bNaeDrUD6kkQtk2mHI5t5vgUEpVL8+0oQfTq7P8
lv1DJFOJOxcrkLFbtrrT3f/YUTI9kbb6I71MOM7GhsdWa+cpuFLfnWg18XY6EoDf+zjdwcVtvglh
TWfAwv7pdqkxGS1Byc7n8D5tUj2AKGLf5rMtGcf1OqxLJlYJJAxavvMRGltYU8nU/yykPPfKwJIG
aMShh81EOhyukzNrUIptsYmzYshAtPTP9VwvYcjR7Scsg6doGChtu0ohg5ftysbzapX2j9MHhzYb
zuuzZzI63RFmpMCmSv/xbfNYg4yoExevRKb1JxdTyyeKZdjDIHN1Zo8AvMJF2SRJCRfl7yTc5v1D
MF7vFmezAFwzwOHTJxqPcXYdBhMqkASEMm4kgggKXZFM0QotthnGSUCehTGxAnlmqnV4A/PODLzE
foDuLyM4qzCSVypllFUa7BWCBh0VZXvbTMGSvloF/FDuV6mrfiNCJ4mby0rhWaWZXTEW3F/cWya8
SPvHo+ozrxgc1AegVZOmGsrIuxdauCdMggj+kHoAxh9E4BYAXUEdGeTi6FLBPLY3KY5xkjgN+OV4
vF8/ZaJcUjue2nhyF+UWdVHGDHY+SyptMFAXpTiyWec0YB1mE7aShy9M+1wQdw+QUfEpee4fPfTG
/MuH69uUvjmYYcQAj5e6MC8hE6smBKPqpoOXN/z7x8ln1h/cWbcoX+stZnVNK8mqF9RJp68onyxo
G/KShT2lWAINE/212oIfOWN91tRIoa0rLFeIPmwqK54PnT6sZOzNVHdX3SlRUcCwq/Fj86Svr0sU
eXY7B8xduAwT1bb/HLN0nrQGCI+8mwWZsl8wVhJvYv2+d3RzUAHWiN2GQHo8+1nN2fTLTnUlyKmk
T76gZGgfeO9pDYH7CahAMv1o6O0TzESUaVMGk42MPdnbuiq9fzd4hYIsLdZiSVqvp6EBuEirVQw1
5hN8PTWbdTbXo/R6SnhC7zOWkah7eqB+YryEffgoZmYHrxiDxFs9vxmHX/wJ1/URqX1H9YSTj+tH
eVBh9yMdsGbWWjfbSTK6bpaBWVNLNKFuT1LXaW2PvXGjkbxZfi82FhE5xFOgJofFLzOTsNSe+YsU
btgjpgvNWddzsvyZ49mWO79YlRgds5lt0Y5cfRUFV6jNbnBDYUVgBCQDWCA0gZIMZD9Mrabv8p7k
TuBmbYY9328ha906ipp94+QHjblcGJfhE/qA0q+c/2JrfHx/jX7ZoCSKbntsUfNe+oGzxqvY4AUi
W+pDmSeGVSG9B616TS2P9Vprz9u7kYZG1GINDp6NKMHck85M1ppdeLC40nUJ72So1bIcLue9BEuv
wYmMwjOHY9ckg+t76o9xAABtB2KDXy/XJjwmRZtqprvBt6BKqJKNSvSOFfkLJv0Mn785q30x69Bv
jeq8dLdnVYZNQdju2ouv4kz7x5sKHzgPo/ha03ffrdnunOab8luFdmeS/A4AdygA+UO8bEFf09EM
SHEw7MttBHy1nI8Rp+Eo8f1ZtFcTdfMnRP9GNMpZVy4BE5op+oqlkiIzOrHfGSKtfAnrWR7cWYzu
Y7G6WxRIqP3keynJfuKYr1Ep+nnOuEIiCz2qjK+lmGn7nmy5ELQZYyQ65pJkZd+LrrTg414Bax04
E6AN0TzBmiXXOpcqB7yCw+zqDhVd3rCQCJhqHjrazLPaLCNA9sBAoHWubzWm6Gr8sqW7f4gHVVVj
TwkWZNtRmuUEZ9BMOeSHSB84gINaMTHoQTMK9tZrpTIaTFeDM83fH/z1FT+QxEzAVfQGsasLuCfG
BYYXrs4HKYK+EOKWSZSU54dSOue3qn3VcOiStAtrwE0PaEE53ltygXTPqQzB3iAGHag6Ef5MpsTs
uScNgMNQBrBn66C0px3minJ1WAsWzrAm+5Wv4QdVM0q7+A7R2i/iumielO+uFSLl1npkwFmVu7AB
Zk1PfzxgVu16irLXnOfS0IYQ/noRjbQ8LvAoHboBmvfmB2jqiomwG833NWV0xUNO2tAWSNIYfp9j
AjyZLoGmP4qsfWgeAC9E6mSM631im14bDt90eok+qFjU+Amfgp//EsMr6MY4teXJf/kfguK7lEV6
hg9K3g3MW/97SAZs3PWt+ibNQyZdM/F7yBum7geplagxlhlOB4Ik1mO2VSmLXB2RdszPSai8q3gS
kCnfP9lrbKK11Od3JVZtJO5U1GRqqnDmWedWflpm+DqMCFClIgf9/1Ns8ZAJEMJogo0XYB70YDPa
6xhcAn+A+vnf8vwEtGjzjRar72ulUaKP99xnV5pblKnQcvqxqs3e1py84NQUIUECvsphKNkruKh4
EjlQeaJFocnD/NhkSnDB4oxjktF4uIneoK82+TTdffAfvcOOJRKzNbKRMCZVdg1Y/FcE8UBke3oO
iezBnkTX/B28N4gHuXBm/4WegSeUrLmEQAanabunXu8a6RRzSzgxArYsUvuesvO2UZ2WFHuZnh4I
KhP+zLQFCaJZlTRbL92xbtZfXR4qTW7yNGC5wss1kyuv5+4TX0Dt7SmDBGjd4wOXdNWnxc0SDIQE
ANwGwNNfJ8U2a21j7f8R54aEOCgDWKGKUibRbhAjDsu7ru0Rup3DR6RgBk20TRNYwnm/NPrNmHvh
HLSYhgGeerpzbmGfUAZztJIvhtYD09wXco4Texj2JpeF+B54jH8e2N/LUvVYoHfrsFiRNEaHkOZl
q4QT7XKrSNnzHkiOrLE8jI01A/OlZLh24X7WfNe0sHYz3uI2wgQMe1GBsOVqNMuvho8isWOYmGmC
T8EKQDlw4D99Z8/ZxlMQYv1Lm2R+drXbTMt1ds66WoXAZcG5EkOgjfJzcTFnAF0Kfm71FQLYm9fX
/HCxONuMVaMtr3xZe0XyUXHibfqt+gx9lyUNmnmuReTj6qBvDAZ4rc73aUXoREThee2nOdV+Da1J
hoNcvSUQ6lEMNCZyp50xr4dW6m7TnIDt6JSgbJDBsOqv21R9KsZ59W2nk01h1mNLtZEhnUyAR2RO
17SRtH/WtMePMZ5SElPA9m60tAHi4yXccCrgU5VErsm2Hn45YJZje+NiLTOemcOe8HuI5FTHqokn
W3icr3pvWcFey9dzhQy6BYcN18Fvoyh6aCbSqkGXWgeDTG4268Gt6fnCE9dz5VI6OxX2nRo5uRnb
7O1KbwWzBT25ND2a8H3n9Y/dXtmAC/o+LQOSXxFWTfDbHvZZgzPMeC3QCj/au0pO3E0mZYgE48IV
z0YyMvb0ApJ7YYO/I1h7NyEXo06Rx2UohfPA6oPkaig0qnwxQuZp4ejNZTSd/C8mVE2MgXL/hr+R
Re6Qf0Bo+naq5blYJG7YFlDjFeXXRAv2B58CIPSe3VLTJSG5JCovQaT/FrqnV4vknswtzGlKjWRR
gS072TXmcLDx72fBpxhLrAWigQorWICjGbKnAMCQ146AmpAGNTKPY8m7dhCS/dFJUNQbJM2wF3WQ
fHtvCUEurkIBCwLsz0d3XHmkL18B4GNAIj/WWt4JrR3IM4wfxqspZxQmadNTpT0s8MYTthtEfc3M
Lo88FeqpCThXlWve1PmehVI6I0NpZ9XWMcNQsrKC4MUqYIHWbv2ArpJXSsjsjtRG1H0vQWi2O2B2
+OZu0SCdBcZkhKjUpYws3njdpUqmQZ/UXJcIQWgU4ImlKERYRyYpN+knqqTmci8xe4SS59+JB5gJ
ksUntOyhL8Z/TDRWo3ZDyFYDqBGkp7Y8IS8tT/a/PRttW4CTf9coS9lN3w5efWxHSWyCTjZWzyDN
7R9CxYrZa98gbg9uuVbwR8xF4bC4FOpW2ljFWgL39qLuFzLAgNu6s4c2VJvD4Dz83Ry8EifucLT0
TcgmswSRIqpyhX1vkwsXEWG55LinL/nX22JfO80jSBxMbi5myBRqM63w8Zg0J78bO5mrSAc6Qytf
8KavXezhTSsPAD7u1ntbN6mv/3icIhkunW9X8uw9o11wgQ+Ra8i8S2GTRNkUOtQJ7j0c6MCCDO0P
c86QXLuG+XMEVoAtaTEoqTT3NluuhqzaZ4F2l6LvGN9pZNXNZdBk1daiAx1CnsVsFryPsNpTt9E/
RgtowcxJLDAy6ia5Dnwt8Ne7X0vD5YgFWtVTuEbfL+phQmzjWMzW9UZpI6GdB4VIg4meKwnFIwTG
h13riiG4PEKgQw6A5YlYsh7KvLp5jSij78fDsxCXmJ/fXFYMxjfNhzXEWc0p9RS+a8LwvQSknFRT
ml4tSHelwrHzw5VN2BkKwkeCHjs4enVM43SGWQDSKv82EsSWHA1F87+RsSyTvVurk0Sx+iqX0MTO
p2JCQ9IrzzH/Sp+ogkKaQzrdga/eu7jve9yCRpoHI2TkhOryGvVrydix/qVuzMTJM5TQIqsnz7eg
Lu673AzrZUi7S6HOAM29KKodDsWhlIufZ7Ik5pFEQmZhfeAIyN3ZEaWYSSQ4sD/tLFiiHbpJFHEv
ck1PT9TsyrdysBkpQX8R6eiukuIbORR0n8PdNrkv83irlogUA4RR20TRcnSByvU/vXVrdPRkiFJy
/dLvt63EtoYk84uiLPg5yVsVgdIn/jzBQsgnDxxuw0G/NTEEZbphsY39xx0VSRcl/iwntmIaygyo
XMM1H2YuyerH4SC/PwsUVfAQgrpNfnUdvXeDlhTKPs4VVRzY5N5KiK8dPb2WMvaKdgiSwtcJyG6e
qjCGNryc5aJFvUT6qn7R077yqLyI7JNQdAVP7xBd3ReEGHJ0wuRJ0DsEqg9dQsnWSPlYQNEDqEXh
V1cyTJpDb6ESlr7NqMEvuuTtQMf1KbSiZ9GnmyzqRD8XNUc+ROIbaOzMwlLd3TZRcFthl3tAynMG
n3yLaMhRZO4a3OJPyq8bZ36GIinXmvcohkFBh865s+nIqYOaKgeb/RL9R+/5Jdmti4V4VmLCJal1
k7Pn5OXX4zNkE1JMmDAVSWStQz2pbotHjdHM0WpzXIpkGx6P41yUMQIQosAyC4TRs3r4qls215Yl
arLerktHMJR9JDnYeKhAuIyazibpgA3Tnr1JCq3kpmNsCD2tli91XiVVStLlrJWcuqSO096sHVVt
DbEFXgo15vUMRZU3aKFsr+9TD4Qf+JVK5Af81lKKwPJb15aWGPuiBJiZB5sHy69qjc5a8PlP7HXC
rgXVJPonhceRNJpDrBQZSJW5MG8iG7fqRUAVcoYeePUVzX61GTNWlZrsCHKWlwbfBnSm482oUrXG
32LnZznG3il8VVXacCXS8rWMf0LotMdxNyy1woYZt9Z8xADD2esAQNurJsmuC+WZSNMaAxujDId2
u0Da3Yep0W42mDt41YdZuzJ6Wx0bqcT7Bmuhga93Bx7Q92LxjB55JIVVz5NdSYg97EiwvNJEdcow
fYSO+e1IZbqd5ze8IW3Cq4CzZvtHcAXqfH2OBGpP8b9hNuQr0gcSENpY1VF6MYcnvzYKCj+0TIOH
er+8ZJ1aR/3/D8PAbwUodf7rl0A7D8SmgS03oeeeVXCZFUtacJ0pGMnoPLC7QHuY5ylJV1wg1kzq
v6ptJB6wyRpoTTMlbJ9qhg9zfZelL5jP3iF2xfzlbs7nmbG9gOiWKPKiSbW11ZLnCOculwBb1sU3
l//1DhGBRrtqfvXcssf0k6sk0mHK5zzVqyt31pL9vjHf0hyBxamkubCQweRu7xRWPeLQKYteQXAH
vklcZfqhoDIcsT4K9YoKIzDkRmvs7q34wWd1Dlb9vX+rQKxOAAlwwgbnDcrV/ut1zhDCbhgl+wSV
wQgEL8+VxC87GJg1vpf+ifCsYAYfhZfJYuKBw7FVUrw4A/jjr9K5Gl5NzQ/ExRomslDhyZFZurEU
UfBpitRBUNxYAZpWwc06fE+r5WxmDH9Dd0wcdZJbWrKNDabpRo60hN/tvHubleJa6TL13g9KqB5I
by+gk3zirIKkMjeileyRGbwcoWg8iGLWeut2rAowSj9ZOVFGcyi+yybET4N+WWSY/b6wNH93HfkP
BzhsICWHoQTJr/2RyCD6g74MFDFgBPJIWErsRwbGv1OujdZCdyeW3k0qWGCj8vhPITFjRVC4Uyc0
Al8KA1HDLWJtJrVaBDRPFlB3aDlyaqDaXppLc6vUne4xqH3Rw/OQ/7Ds/XaFgJIoqt4ZmJUVmqeL
9qUijNf5o0Ao4l/M8Ta0ZUi863DZOGG3DKp7xNc6+X/IT9qlVGqzOjfL1nzVd/4i0f8YAISXhsz7
o9ile1QNjvJ86hdBzZcZUDtdD2AsymIxYrLpK8FkU3x6jgrH8Zll7cVmYhlfRslSgUYadr9/qBRt
kKL/OZdD6eHwtG5+cLG2GqdzMJlEV/jVmYU5Xqz504ng5zrL1jUhzLSW5j+4LqZhy0zdQjsO6QqS
sWBTaPpof+7spVAnjWyo+5ns2IuW3y4XrMqTR1rZvfqfCgp8TAZ7/JsFlpUT+Wfz7qgcNiryPvi5
nva5o1EwFmHIVGtYP4InLM/wdmmGotgc/bKpL34szrgM7N5ZJ+6Fa0BBXs7Qfab5m5bfL7xARUmy
aACNkXTO2HNG4ZjlMZH5BiiEdDAAmQxd8yQ2LP6TNB1B/abpMgIdggnPsQ2Whwld70VpRU1MVTFF
6yYL4v73TeN8wb4v7GK6jcw2xuaPtlxpJBCnFn88xwOjwh61htGPWxiVs2VE6rJLcUyx04Ci22EE
zVLkDJ6zbv1xNGpy10VRO4527KSSigWt6rAoQTHI2OlE1Tlyg2OzVuu5iy/L/j6enJgUoXXnsF7b
ezrRXDmPXezIIC5g2iL8nEFMmXeldNnpeMIuMez4S0NNd4G6ISMO3gpZYeiGWjsU/pX7DyTLTeSd
aPOF//blXwJrOfu9vfU45zmdnFgA1hCGsk3E/iXnaFSXfqTWFOBA4lieUcYRujRfG+4S8JJgaYFo
UQO1dtrzbVjQpzriisFPRD8R0HDHCnysqhwb/WuMl9fMFaTw/NhF2VVbEAqQZfKJsiyY9+4GvxIN
1bkpH8H7q3QZlEzjGEET8M8pz5tlDqNQLUQ18BBFh01nuCy+fsi5QY+o1EF7Tt2Tccih+P47/jMt
HCPBSwaPBZXpRo8VGFiSqlPlbDdwR4q3a8lVFVHbNm9t6W1Or2cH0FZyWGT+peFabQ2QGwxdaw/7
rXcarSyy3bS1KkMM8w4UON36MB4VYpXFp0NV019v1lUBcUlp291Io0RBvKI38HfeHhgXCOPE0D7A
Oa6WP89awwnKsIVgaCpHYi6wOnD78tqe2WJgyPuD0C4gw22QALGwiz/p2938hEa7tPbiewBafw34
6LUc+65xFhmr7bhTYkKsGhjZS5leuz7SUqbqR2xBpB2PZQ74Cv/hl/WMm7Wq1B1YSgKSzAW9NGX0
WF+5wIecx4QLmO8mI15y4Mly4yC4oZg0vTOma1n1S0oqmudoMTvvlJe00SIoD9zoJBpRsKunFqxh
+E4P2rjyv/H4PJJDkOi2G4Q07qH6bfue0gkpKkfle0iK6VZRBUw0ImJ/t3ZMcvbtObPKvNZGES7r
H4y/nE387m96zjI0zj3kFiFri3jhmnW9SxgGbG5TZpkllZbBoHFjuZMrB/s9CmxDNm20ZWXDPLa5
tACpbNCC5+SG1WjGlmscrfZmkrEOuJ+FJ4LWz6qTwhRdbjC8I/T+JkuAbZalxmw9wimt/WqDCBZs
LDtS4ajo71nRmfjGjWQA7ZadX095yj0p6Cvh7aTUB1YLfPAqXMmf8/Iu7cLyZrKC4MOCjLjtX0FT
ZW343nif43DKivfFcsAQWCnS0HcDFqJCcP/46ORhSCI53DtMZj4mGenubJkLqVDmM4GA3VoMwpfc
cwsU7P4Hl0ou9X+uYxGLj7P7T2da9xk/B4QI2MG5MPJ9hS193ILXWnaA3MQdgyA5XiLp0PYk99zh
Aip8grLSkhLrFdd7iYpk3hh+LzLqdF/F7wl+wH/Cw3tFuXXrGGII6rWwobmSKrHV5qtsupCADLp8
MSEW8/gPydIF7UbVJ2rcOwRPxpDpLm2c1R/rlZShF/AA0l1HfMKYXsu5dy67rqnLoTTnvvIzCjJo
o25Nd9mYYolig2xUm5Pmzap+vofY72bQKjpWM7hpwM1NcPYdNVC6PJdWTtoXnknm6MMJI+SvTgBS
bSRt50oiqcSlh4zwV/pVH3pNChKakucywd+vbDdmLaqGkZxYA5lMHbOGzq2p2exShWsHl6O0EcHR
glk2EhZVz1376SFRsYJfqfcpUppyHzTB+sDkDHnwpr1Qb4zA9njHebOIO/VOojVvNPUn4mtJqdRV
32qRaqfw2XXSQ9bsLEcNWe0sWRyESpyhJG9jMwTBIeoE9JbJ7P1cqVzD8vDNrnINCZGhj7Ux03wk
vK6uV0khT5ZD1zGDIOeAw781ruYm25kOVKJ9EO2A4OlNKwC3KWhcw3w11j7a9s5AwuWqRgkuj/A9
d5NC20jx68axFUlocv//sRFzdvyrV0ii0tMxy7RP5DJ3M4xtz1332SZ6rfpwlp3o3PyZ8zJR2jzs
/1cGHjxY+/z3LR9V5T2L0GygGf2SqvvjWYyCTGTzisL1obScjwLVUdMWrbNCqCxergLqYOdTPF9P
veK3x883JJKyX1TzrJ7nQiVJqQzBQfnBmRrEIoai3CSPXHk/iORyDNY7ioGwTwpfFJgfvcfFb2MP
l0zbc7XB5EDPMT23IWuaP+oubMGx1Ir5xiDqLsix2v1+x2uI/eqhb7lECM5NbbsxfsOb2K4/iVwz
+cMPW7OTtXaFHa3e9yoGvj2AouvPkKUqe1+cN+ag6h7GsqQ8Z5p+Jl5PbbQcPcvAIXhVGUc+t4ps
0DwddHLCyN8TF80B6vC56AHD3u5gza+UOr6G4qor/6arj8j9fpQ8HOQFnNrS2ICYibLRjyHYCH7V
TwyVAaQEvZCYYGIyTmlIC6Bk7KMQC9umG8/BFJ+z6PcJzVZYH7YjyDAa8q0+B20EIeV8zSKXfBdv
+NLGD0F1lbLkhRsKPOAkEgxapJBZTl1hrs+UzxHQ6ulO3LwCP7x4SgwtV7qhtNC96jdXHd7h7cQg
1aek3BuMQALq4+ts2YY4BCq3jdNl8s1rnKublLvLdR+WM01qqAGvRaCfI5IybqFOsSseucZYvXKK
9Mvg3EFUUEqs/axMbp4DfL0APulRhBt9U4kR/ORgfowJSqySwUsG6FC/d9VrmOIP51/nmh3ZOlMB
06Au5WvFJaOGiphK6V2y+EIqK7Kmwr5xydJwwM5IHJZ9svlqJw1t4X8CTSUAFUnQLHerDP/3928G
lDeaPHLfX7MhnHgX0ZrbUlUGcY56C4J2JyhFBbtZ0D2GaEbbuq3brD7yAPl7ji7rA3EMMZ4O4wPZ
xZW0zL5rm/Og0Xcz+enHwQuBQ7g0ldZy52cYq4cxsBOP6G4HOZuHl4WKUa7G0zeJQ/C6cWYjkaS7
3+KLAZOy53Rg75YP14XM6WOedtpE8uDf65vUK5wiCAlOErhUAPn9RQY0kwIeOTf5U2rpdztIHNLr
4NvcmEsJiz/tbMndMei4se4cW2GHaSmIS68SgK6gM2/i1/Z5W9ja7SuuVSiCUEjgu6l6lmmC4Hts
lDac2emWpfDzNR//3dXI81DX+1Oa2v/TX5vyv0y1ju3hQ67Wi0wxR5VedXL3BMhWTQm/oz5qZ4u3
JeoQgMBaiRQsXlEIaGHfVcWjpvU5uDRyTXC+Ote+THHPbdlONOGpzx5wT73sqY+aGIxZ7m1FvrK0
5MX6PJ+gB1nMnR7x43LENAbq+9r8ZEsH/DplOEsTTg0P7H6rfnir70MHDt2SvDeAiVVx4MQuUsGG
hP0NTNxaPdbIe7AKbO9Y0RFyqo5B+LXlFqI/hpIT/dB8eJWnR080JdvUhei0NbqqMM5/d++vAY8T
xn5AWR+6xGzI0ednDEcJNXFduOUFtaxD/SPl3xSdCxwZPJkMHHm6Xa66isGeE580vTT7pFmgBbDr
aUDWnFazaC15XVK8OEmu55HfyTAfa52Vh/PgLTeMJCgLfZVRMP8qc26ZjX+N69aKncFAhLE48Jal
02QdT1YoJMh1M128KTJjphpElJtCD2aygRG1eX/wv38qmKbxSkbMfGhV3mOoiWbo054kRvYbY/Sl
FdIzQ3VrtxAd2AguQdSyJm2dbPkIJ/LWXPxddHfYEHVzUSih4m2r3IXbZKaY4ECpKksV5U9Zx/ij
4KcgOIE75RkmprZMJ724rlFgTtUfo1nGpnNsiyjigWYPPv8ekiwT3y59b+1pelZT7CncquoYiQUh
x2m9j3RLpClFE+7DmAyy9k/zpycmKnKp56LrGkev59HisPQFSvQNAqf60zNbnxHy3xiDvmA92Rrb
sM9gcBOrnRygAjU0jexYM9hEVBttxfCxZCQn16+rqyt2RimkWWlBk7CIxhcqpQF6X1jnFiDaCJvQ
ON9mUfyvPD4WLAK6a2DOwykpOdUa5kUYXWG464vkaLPoz6f+3q+V8hnAhg4m4NGh/20d39RIT/km
FHl9aSPMDJ5xl4eQgyk84db2iXcdSbmVUKSkvkvWfqNRHrzTiykENyb4o8o3ki1MB9fUg9XohEUC
OiXKoVoq4pZczvC+mkXcufbwdwbBit5Ca3QnIM7hjU7k3s8Y6VHwZkxnA/PFUNqEnTC4vFIf8ylu
9FblsnGJ0C5R4fxmGOlhqFYgh4tiFGJNe0JFqYxkLlb2+DwnpJ2xNLXCvQNflpem+MDeNe99q2wk
xEfvOSKD/J9qmstFhRzJubdPWtnPbQnJxQ7yz43sxt+deDTGl5h073Mh3r2qkG5EIdpHcS2E0oPY
fgXWokcecvOaneDj6H3MsQVjkSCrz9+Nk/OScwGuOTxIFkvcIF1cL1HixOYYIyUm9Ms+gv7yzx82
WiODuIvwiVpFEzEPbtfFuqU58CTkj0BpJw5YK4xz+nZlJU44E4rwPPOxRq01gperadil0w9lifCE
YnKyI1vWhZ8baAmCh8FqQKEAZd4YEpr7ALXZuVbteyVoK+vcYAEddST23iekKYHIxaQU2p2lNO7w
6vPZ2x02qi4y924/tpG6waJ0eyZ6Y4EtIKv6fbzsDOofv1+WeBlOr/KEP7FMiQcUJHAXjDuOMpN5
txAk5QrD7hq4VLqqDFoE7HvQFPzQD+Aty3OH+zTU9CHeG7/KnYKBpgOtZpfPIRiyP5PP6lsMPdcK
DnA308HF2Hf5OEPMeUIit5uLAvRIUmNGkJk4QHfHKNELq6pkeN9xzA0ZtUvz8t21Hq75YtInRAiR
KqN6SLO7vLM7Xq4QYR54Aid6gTBvoB66EI06Ycm062nyqGWiS3/jPV8CRHx8f25Bxbw43uYlZ+9F
yLneXydMIlpVFlyrZBLnLrwNxDgAKjJ1uZym4DmVnSAwWLZjONLBD0tnjS3WV/l/H7hU+HciyZ7k
6+1jrc8Jk5QPnNH7SyxLsAKQe3iBO8Kmlj/zM/ehHw7pAenz6QK7hLLAx1eOjTs/F/1jfjOdGKXL
ksXhDvm3qccRXBZ3/Ju7YA9UniKmV4qrq9i5IejhXasocF3RBbvc3D/fs4d7Y2u3zHANXiz28SII
6RFYkz+fOLUx4LUFM/cfGKbp+pI9im1lxufINy3RcdWeOnqAZUOUJshkeeLnynZ3DaQyaCnXm0vc
0NJgI5sUPdrqsONHXuUsq8KZA/dUnFSLNtjmB248dPNS8oaEwccayxRnOum7UpjuDBnm46S7H3yV
8q3mWnhRKVKp8r1cKVHMC5+zfvxCX3S8MJRlw1IgtUTAFDWHDHMgk73H7rb7pYuJJYa7SvrKv5H7
5eLv9kgd5ta6FY+4DYX/jUdkksSl9lfETns56PIGiLmExSdcLBc8hsVwiRBdgyt5zBC+TCoaQiZb
lDCiWU9O1lUkuWSm4QMvPTusBSaphBEwwkYb/mSg0RtJbX7IfyE4gPuP+7yv2wyNa+g+cKX1bBUm
2NNd/+VUxWJmivcmRHvYh03ve23av28AyeeUxlnRViw4QL45HfmReUBGkJ6ClfiVhUVnQr980ljE
vG6J7aMo4KoD21UnWZWFiR3mRJceSu+IvLEk7IbXkXQW9SaNfvhe00S3wNQMkmxxS5xjAVoW6CNw
Uqf9sytbrFyP3Jps0x5tUkXk+qQxFEid3CZvwBqCGRichKIDdAowy+UH35ckcAKO7N1rGGFtqTf/
kT503gCQC0RgEuxgLqFg61B+yOuJ3cnownH9hQvrDbr3CpUZsUPze+SgYsHhCQ2LqsxJiVZwJACQ
JfB1oS14XTCx+g9PZuGP5HBY6zuCuv6xufFrRjt0NsKIpeB4YWgH7O2jWTLQF/mY9UyDwrpfPkYU
9qr439h3xkH/4cpi8XOlL+E244p0pwhSK8/wYk7gE+1dYNWem3keJGKcdrQxePD67iJidF9pxOFC
gWf5+h/BtRWVWd3WnLYxWwweZ8iYcxEazR7ScWktGyJh134YoNQ2yxu1PS4OurGAjSMoL2hjkC/R
Ubps1errJ6HVBiunYHrOEmRA93JfPjNPZev2tI505k2cC82zKQOm9jEp0m2kQ8GdToQgD3HFTRMh
N5bFQKW5M8ms5rRJYVEl68EofCgEG/EvJicVHz8//w17NhmmWvzqibuKlSYSwuPb+YgkBS9WvVx0
mn7Yp0MNhC1WXM/3wY40EENvnZj+5E/ewvTIpGRnkgei7OOhXyrQinK+UhL9PhgabVBeQgtpDrLV
W/XLRPiAju1BmFTFPU+1D8nKOUNQMnSYDPFhEtupsdv7uilKWz2IkSq6GjBcnqZStx6jn2PwftfS
htA3hitYbfeLFz+dLpjFO7EPVV9Rzl1ZM30vbxqv2ZQwo1Q8kzCoHIWap5iooVaMDHz1+tj3KLAM
6uM5mg7nrjt+C/S44tUM2J8XnPi9s+xg2UorHcrj/2xss6In+0SPeFLkLdDLymFNYCagPjJsZ6Ig
540F0ur/wszM+Sy6f8ZorRhyU5azfdo8hegl0Q5GaSORRKlpw7aznSppnM6J4hrcg5BsgAErov6e
zFkl1fTccsGpS2pJ8smEMTFsjSP0Vu2T2kDpUCsShdUCnV/C+PY/CF+eVtEbUcX0siTPPPTQqdBO
4yjwmHfSHIocYB3QdwymlX+qiNMQkk6Y3zHUgLjRhzh16SfdvgbwsrjF5WxPP70AUJ6F4ENZIXrX
NgfNtgd7yT1KO1I2yECkhl5NRZ+EN6NgBK1mHTbqzR9FDJHibIOKvtb+KJFT7st1LQ66Mg3CRCxG
CzvBf3Uecoy7mouGJTHCAvmlaaX7E7hK37XVC0jzzBRkRqzpGcgRzh0zO5Il/WI34DnEyZb9xSlE
8TzKUK3B9ZPGM57UlIjr52k8iyqdhmYIzrTSYDy7jbcFvPoXdDWcfTIssQ4jxygudSft0W1xswki
HjPLea5R/k8SONVQ4lK7lCe7hFWiEhqj3XDw4qunRQ78J2IVsXGvkaKw6Rob8Y02P836rBkTiLFX
Qj9u3wfcYn9PJUrarRs0CXBi2uf15jPCD9HPKEKMzA1Au9KVmhlJ3Dn7DcEMJJOx6s8Z7XWuYsVi
8SkpN43m+bDGKt2NJK3wa7nxSecJ8Jfcd4SAhUqgsJ20zURA+/OeqGQE1H0wfhI5P6StoCZ/YZG6
Z//5lOqEf4PoN9Gw/Nw/rYgfjzzhXXrLoLV9eDBbeuyFsQ3gm6lWKZ29cptAJP0drkpkzb72zTFD
Eu/PEEp24yv3QZOyunG7mh4Ec774nPnEn3TEz2E7mDi6v+8KTmPLJVnBEvU5GO3oIYr6DNwwmBQ5
g5nj/nLdyV93IZIboGB3kQRXCLXc9xzEEZ+IveDLnrxZ9Q3PDcMoEx3MfpyDvJIiGCmmAFh2oQrM
6XL7HScYWfDjW4w6MT2vEh7saZeT3UBdXrYcXbMg2UjFvv42ok9bA+C4A1RCGkfCixlmE9re5ZGU
svqZOFq7fqlNlvuB/M08lsAzXZXP7Su5ntJdn3e0U/hq+EbjsMpcewEtLtyhwUTpoDgEreg3j77t
55fABQM9KXn2oCppbxluyp7CXhrt/QwKSo/JST6rabJ2OE6bYrT25g64jYYOKD7fB1h+FXCWKsZK
+7ZZBMPQtKnh0HqP+ST0ii/J3ZtDqOwcYgxAM4W7qghm32/mCYzNmnjYHZhnEHfUBmER7qnZ1V2z
BzChEESM9T7CUToJAhYzePAldKme5XWMAdL5RuFZ7dE0lq31YtZCggLDgfhXAJ3hDBlh9kHxiG2F
4BgutFqYLgAfXzBanvTHKhknXjD82CKAlua/LXX6Q/ydMasEZTpmmWNLO2JDFMiMrpXmHbOot2Qm
1QuAJcOIdPdn+bLCBfDH/Z4eq6qc7nVEkoU79ztpHjccRI7c3C+nuiP4cpmACXyLxf6KaPkQ8N2r
jNGjluaidmA2/1eMlxN2AsoBzrebt0sKitpPf9Y1u4cK+y5nv4aDvLTNGmWFFCzkvySO1k3v/qUN
Pcj2ce7If9fulocSg9r763RohgjGmnEouYM23ehUZt6QwPmI++CQUwXZdL+NUYRgkuUmVchYp0FW
4HNSjGR7EpIeaLr6yTMgx7Hjb7VJ97/UdOyI3aSCXilkiPe8yTMZ43nXzRAboy0133Ie5goDP14P
mPR79nIqlljC/ltywhScdLlJoCx2DKr/QRhWxBi1rD0sBmr04FyNiMfhAf0SDf5iL8xgTNYakrZJ
Xun6hYihwL628DgeezMhgCigrdMaQJ1MJRF1NfCyuFMSgf6EIph3JsG+3KAcHLvlwyIU9ZndDf8u
J2W1dtHPfwybpcumEz9vdcGGvW8rWdPxosbdL1eZ7cwdLvDX0ZA+WYq51tdKcQwOD12GsCjHt05a
3JcUrDtTLyKScGpdnhkmvBFEA8s1oaI254KEI/IyY+RpxU6kQ12N5oZhlzTtG8kRKGesJdw7AMlu
Byourm9GMPY+gSdWvjx/WJrYzh++AN+nU1/1VPCZ6zoScGEvdIPSKVWt7mBd/Iuz07pP270XspRE
R+GLJ4CHSyl++090+YnFj+PXaqcqcj5nU/3xNTfS+7Sds2QY9dpbufpOfVBVNzlYzLS8EOMC4FYy
jIji5hDWBwHWKJ/eBSjdvcBgNuAeujIkPvSpEDxfSqRGukIfwF8WDgMZrN1prd04pgNQD01ZbQR6
r1sxkRXg7SxEHWTzZUt8/wGOarA3yFnDp4mBPb5psfCQ6xUe+eOo4/eYG7Vl6Cyt3InsOddLjcAr
pmY62vIM05z/hHfV6q7PPVy9+P6g8BJ1GckDRosEEfgyg3f+EKPejX68c6eZYm+isLakWHwp3DRF
V0Onb0qLv3xRjJC3J7nVdc0/dV+Ciha5xaNfF3T/o0u7ARzZ2P1gD2h243R/7dAVJnXTCQbi7Qg7
iL9inrfe2ysIOhUqInqUynup9DCKSh9YBXKTCyHwxItlHjG/1Fxv7lTifBqU1EMwSyKywRibKuaa
/KsC3X0Er8A0cDjUzhIJq/kb+z4t25uNfynaIwLPusmKOGwPMIS26g61YgdP7KuhSLPbAL4Vt53L
Spz2GtjhVeCjQAqrwOnwkQ2Y6xtEEC2jVsB4aN7Fnp1u2h1xNntscEYImuuHc6S1HA9nGjGfmFow
i09I+5tpC/Bhzs0XSyE+jPrucQQR40AsvL+saoiLf2vs/+dWyCS+QhyX4Becju2vFODccHYdnVCc
h3VnZ3UTx64o1P40ZcIOyDGIM999HAoLr3fHsbni3h1VWZxUBggh7iWrrX5iMBeEhLhECb0XDRS8
wv8Pnvs3S8DGCgEhc9ZWlqc5e9aYHFP5KE5e/0Pc726NSiFHpFhCGWA/XDcB3pOZzowsvdWplQo8
/MzTSoqoSkyZ/I4lvFLnh+vGiuEegwfYXmQ61pfrI/1DnOUhw0L1cApOcMcCmYiuKqSJF+fvmlvU
trUVWwSeANpNr8ZT9NcIKARluEO4I0q9tF3B5iqoneE1ZaX0dxhmd0uZCgxIzTMxpznAffdfbOhM
aBRiqDNPAI+XvmuKi2qt9wx0AErML4bf1ChlHimqUl0VigNunyZkVh9HzX+ZJ6Lw6J1MHKXNECMC
SbGiY7/QdUu5g5cTnjcmY3YrmPKLOPRtZD4UdolyN79mdYD1jjdH9tgCS2yzTy7hNtHCPjYdNwlr
paaWWRLv6dpzPjMKz0WXMI5DeAW6v3b+QyHP2lrolqgZhEROG+iwxYOIxetr4JUTf0PFa9hupXeN
6Q5AYIrteiylKJ+SJGtZ+LlGKmW9Yrjq9Rr4uMisBAHyJfX1HByKh7w7wRfd/IarlhI80Swu66pM
mgRAwM1FKDzJuX2yAAT4ISriJJI3tlQ38bgw6kVlnE6gRE+vJX490nlN/hQS7rpWfjz7SdA0hWS/
sfkdC+vi5cUUsSmw5WN5tE2tH3ILDcnhwoA9cu+Rf0cHSPdKKvRgzHRSxb+9Oyr39DFH67fhrdJf
fKLDUyCoE/annlYVUf3bNNrWdL9SwrkCt5CVYome4WiTN86ltWI8XNEt7Q2Zx1cDx92DsaG3XmSl
v8E0sFZ5Z84Ht2OBTgjEd3d2k9ECBCu83TuJ7VgCr6A9GAq045lwh/xWcoLbtS82KCXP33Smth6G
Yw7+0sVGtxTrjJSuxJ5givzgO7Jy7bB2IVudiDiXI2sB+kA+I3KiJmLEzJy8PYCkU8QWJwmh6hiu
Bbd0bvlbansRSYrX3KmedslHmCP6RtYkVFc1rWLk3A/4Pq2OSGzAz0WFBjIJ0CS6BKZi2hk3KC3j
ZcwWzUO9xqFRtcZp3brbzeWRlb0c9hlZdGZ9Tx92mHH7yvsrtxYkUMynIg/RqmiQCC6xYoi0d6SU
x1nTqAuDZxy4mMtMzw8sdL6tJtWXd/Zghy+IlqH4vHSvDxPNz/XxnLAn1Inq6Q/VLz02M/iMIWaj
Jugs4qa8KJ2NSql5uquI+DAON8ITNK2nE9MPK3rR2LeQogIwPYEipZSSPqC5GixduhMvB1g4IWHR
EiP5gzg/J6zeh3HSfwhUXkED5EXIco8hKGVGNANRLLajNy0a02It0FD4iYaI/KryHb4f6uoxSX8A
y189x/EpgVEEF/As7S+gNNxhMVBqm/zSP7J8LZxkGqRyuGjWWLZdi80nAnDtm66xknEnunN+5BBn
OXEIvyZ+IxA3C2tLqdjOl9EGLiN7vDil9K4U8csKk8TW1YxcMbNisH191ytQ8GhzxTVoBho0LiTo
+qR7m+a6oaYyHGB0RBEEp8l41vkZr//9m+P7IKwDx6+LV3fAFoscMh7bUYvy++jHCV5iVjQpSd+0
ByluOKC/VpIfbTKgmJFc87w028pfXmcx3B1r1oiDYkjE4XjsmSTFMtWpO1UNCZJhKLWwEm6xzAFo
y5YGFmHNEr+RrbPsBI4cz8pnB9+FqFAt7io1MjleGO/9iZjj19YURKjP16pAOtu0MNrQXsIPabhW
eljYRDd+2vlsCjPQtyyKddHgwm3C2wIJE91inrI/bgMl+bqY29eHc0qXwhJOuY/2iPmEOUB2zdNQ
+Ps0xA0Yf2N7t1w7p1pty7gKKuSdxHp4+2COotODQIqg/NDaa3hUATJGEGZ+1bEXVrK0I8nLqoZ0
Xh3feRNam0Ip6b9Vb2tXdL34b45sy+5Pm0RzSq0vH0qpgEr9WRvNeA/masOpuGEPprFcT3LKSZIj
VEqJnBBiPkofUtiZ150F8VjXp3PqNlQ/TNA/iVaIRwuGFd2sK9kN3T+7XfA1Xx+BZOOCx9cn4nTv
YKeEUr3If1TM3iR7BYr3wFxaVgewIPR31MrmS7pWX48XF4UybjRb3eUSg/K0iPl7re4RD8mJwx1/
MA1bPLNz127fLhSR5aX9nHYjVRzbv7Y9ck21ztD2W/EtRID935ohek6aMHoAEpRIQsNAhPZwyFYU
htHdH+a2GyXONVgS1n9/zFa6wMI743Z4ikje4NU3DTRGCcYKOr7w7vAJkABj07gnFfQG6TutgWio
P5MTy8KOjGcatJwzvqq+iDAczsM3NufBx7A/jIiL+tdeS6uhNN/2Jj369yxsd15Q3hes9vPSyoGX
IH0ZRDV+vWvFda2NUyx6cBCDL6QRMJ4OTKR59VQiPG64mXu9q3fHzOulQNCVZQgD9Fbewz/oTOM9
TYmKgHc7vxFCkuQAd3LX+1JhEQoRtTzYkrI0MOT5hzFjPGGGXXzULQpwdJwz7nTqzOCQa1XOorie
5CMEOFsBzDA/M/GaocQYpcV4MlZRzRndoIhQMZJcoVSziEBV2jRcPF3+Mrbbs0fjWPEqIBi2ZVuV
t00oP5+fpUtyNW/TQ6SJ0oXzSKYyUmo3CQ8Jgpm8fWSAhZSRVvM/pT8j8fDdquOIvZlz/8tnGNPq
BzMu28+NdDSSrtKA4EwUfnNwwvn2uIPqhFSuDm3143r2d1cYhJLt8c3xP7PZhEHL+alJPkUuATLd
o/mhqrShoy2M27cUX6PDEPhaUzyv901VRGoF7JDsqqTOikJhK2vB5fxTLctUwjYHphAoP9rPOemf
XW7kCB07dqK/5Dfuzemzu/6PEiIttsPgrKj0wxYNPItOA4R8JdwrA0Eawsjfwxu2a7c1NEqDnR6G
iEHP0Z00zRP/r5pv19GCYdQBB+lr5XG6MJn+jXzamnA/ZQbl7szU13R8iT84Mjdl/MM/6iWWg9eZ
HmeUfuG2vD8d7PtG4hMoO2xmBFwZwnKJtZeeFMyqz/P8xPSE/RKmzz9nED9GiMQT09laF/vx7cIX
hP3qooZZAq8c1zYRtJaLEn2GdEG6Af0rEj3mADDB8OV7N1LJ23xLDLLcB5RCeBllv/fb+PxaIeGk
+45WMAJj4l4tGm51u26jaOKtk96WwHOQxZDhRziYwjQ4bdPtQIrS9A90C04j4h3cd33ehBtwhwlR
lUpFZXYX/WvV4I827/KscdYT/21QQoxmZoIrs53hbFFBwJCGXv9LSiqTa0VT7UVIsdDZ71mfhoX7
qL2/iVcrwR5r4U30pX0itcQRWg9hzVKWpIWi1Ki6U0E+fNDl8jOgFzJA/xuZA2EPh7o1NF4ilFd2
Y06Ps/YNTPBVnsa3XOQmKQtyfoNvRfldQuCgjefG8CFOx/dbtIQcLM1ajnLJljex9SxRV1RGhKON
ckAJxAU5cVhmg66JMyy7oJNIMZ2FcS00y6uyymUx3fZqfO0Wg9wVCXHmvMVhoAifzQ8GYP/lyw9f
aBaZTLePd16Z+mOntCpvjBIGVT22VqCxBSPVUURz4L4CN7HttS7oOToMbZtfg+zDdSnBgBY5AAkX
bN+vSvdLIgXQVIAWM3ILpirJWW4dCZxIXKonm4rQ4335X8MuG4SXip4LItveG9PebxUVOLo87lai
fRAZkQ7mEEAM5hAohSq1G0AYm67MzqI1QDgSxpj7ddUE2G7vajdLPPSwr1xQqVTVmXRpJ3cyCUa1
2w2fM8ISzYFkL71mgks7OHwhz39LuIkUU5mseZI50SlRVzFTKhO0NEU3mWE6Z5FaGQ2ygjHFxTz3
vQqmphuA1+gEoMRX7WJQDlBZhjclthoRrOxrvAEnl1vn4Z/1T7fEE/F465rao5ZSaRAcXqjqTLBc
NuLq9Gsf/YQlzMNOlzL+nzdsgoC3XCgpM/n6AJ/WS43k+oBkJJuNTSrTdutu0fJ9nQ13iohu2uqT
w5PGX5zrkUbciqgUDHloY7RDySpVXDE98+zM4uJmkpL1PiT5b1g7C0QVXI7LUgCfHTgzhigs02a6
/z28O42QCZjZperaemmRcXMEwGxroZxxt2xlUKKk5K/P/f8vVNPIm2vjWUxxO2taYILFJs8NQdUO
Su7d1JdMn6QjgDA2vdioWKIuer/UZFPWOye5LvM8uEzFAKHVFdESiOrf8c+P8Um3GnCRsbZhGRlA
ePSa2FhHXdicVWrPaKKhNU2xQ6IizIUi40Oe86kteKmHdnsGn00QloHrdLUPZOIv/wOUNV/uYwKp
CQX5UKMtB3j2USyhJmVG8i5pyXCHMWXDTk39BSrENH1yTYsLBjH7YpoheLyffSAfuR28X5WMZAMU
fnd/CVic/zL2WbcHecLO9x4LZvFjnSAJiDeNPcv/Sfst4z4DT3fQXyftxGizJfKdDiRmlIeRkPZu
6wyG2ii4l+k8LDy9Dv6ofEGjVxe6b225YrbmiYd2y+bCJMHHK1UUIWhyodsbyf360LWtOGApU+kr
RZvncfD0I1Y3QS6laVTDZoMWjPERGLXUrAbXgGaawDVUBc7M1ObhQzdQ1fLIMBXdZorwBjdx5fXD
1nkIcVc7C68vjgnhBGgBsiR4LIcQbGlzSfHXPryBFCR/cDk9o/AfR7+sjLqTc3Wa2d35h/S1lpmX
Cp6eb0khUbw5zxVD7bLj3gqHFK0j6SRRusE/Z27oQosOK4rJuO0hjYsIV+KeN8mFuG/G/QH+Z/+i
bihJZDPggXSA0VIarCD/VSBw5p3XnVwFwZZ/E+RFAPV580bpuFZDqc5nrB6OV+abpxknCkkqbbNM
lj80lGL3yHSjIL+32ud+VZkaw7fpPzIForhpHEqRf2FJ9w8ho3G2pt3caflKUkyr0QFdf9Sa8vGe
cC+tfpJ9Sx2T2J5560D33s96tC7G37g09KLacFKdkNFoSNyf4kGnYEvzQCzczADLQCHWyTPCrjSC
nOGRbaiE0NeDgQc+TykzTw/0nlIHiAm+nD5ww/FSNCB5vI6BppJXCz1ayvV90nHnVDEGg+PA0pZW
DLlisiSn4wLhQFVTiO7VooVB0qYF5WQIDSEoihLuzPhTAllkgisUIbZForL6pC0kbPbZSJK222pI
pcy4lMdxiL3lF/SwXZ95ZJd3X6soJkRrPrG//IbFgrKma6RSyEZ6w3Q+E+JN1Da3dTQ81yznlvNy
MrwlWX6COzbMD2awlX9VSz+mVm+d++imOHDcIIVVFAy9vb/LJTDgZE7EDumOD26+N0NEKjR2MEND
yDcOiFqfqIAG2T5V6KWF+bb0ji8wFkDhO8OdLCm8gI+rxfxtEZwarJMcQTHsojnh6TvO6saVCvKH
uhc+pUPaofGkqd9/Qiw9DX40KmS+W5rfs79iwMXIzCCkRJKX8vC7m8hZGfp3rh2ia4OHNRvN4FDj
1sEMW3ng6AuHWFW7Y9/eSIkbNEHucUEH4oXTz6l6k8Ufz22hpOpJNhyPBr4ZlhcIo6Qm8UiI9AEB
hOc8RnSiBqS3OuKHlYUjDsB6sbp92rmHfaqEzT3+B4C501ZrJhMTu4ZBSST5nNmyrYz65ExI9p7j
CMBQ99vqtpnKBmxoc+nM0uzuh/VYZSivJhFHA0cMrogYIaFPJmo+fvxkKRmhxbF/zrBoroTkLWXc
iGsyPajqFgvfEcVTj7AevNuW7OCn1NKi7QXtXmoJJxNk+YHOhWHG96978ffi3HO7IGzoa3fQGG1Z
e9xoherMu5f4d5VG4hcL2hAQ9iybI0IxWFcbEYbMzkeRsDU8m+zkMq3zrcTbCZ6+iHvzCOd80pvE
C/HIieace+749qi/rRXrw4FKTn3Cs9n+M4m6wKX9BNPqnx3s4GFhkL0/e4xr/j2yNyVXl0iGZx5j
djkxQ90pq6u5dasp3+t1AYItweC+zHYNpSJMQ3cZqDRQ31vc1GU75uOjUlCnqDM8IYvItvjHo140
GaAEbm9sTwUSHlDmBIF9WaUrxVWslOwbdeK65mGQ7UCpXFLrxC7rVUGp5zsX+VQtpkRio+kutwbV
wgpzVisFQPpqalGuIT4I6FN1iVx+5Aq/1h7b1a7sG3KDDaodX59fXDy+UFJGD7FbS6CmTLOoliOO
N0yo8ckMrksQeb/b630gcZ+204JbHvE7XKapkCZoyRQf9n691Qe6b1K6ID6tEROwoVpSfdTAq2IL
JrzuHcMU41ehBEOaKbkX0kBlPEk797uuBrSLwCNGBsmgnieMdqDPPSq369VZuNW6SWukTpK1XGoS
3G4uta8dkvNqdrV6FUMZE6NXRdvnx0FuJL1M4go3WYYDO9+tcwKsrk16r8Mma1eHfka9LjELuikM
dwrXhBfwkhH7oNJX643hxezX/6dguZl5GzYiUm3fG9BN5dPR8xtSxuKnzlzv9XYtBx1eFIvh0P+9
BBaTY1Ww4yM1dGzQOsE4pxJ8NoZC94u4KyuULxaQxOxku2slE3ykPOBGG4vysaXb/t837icq8pCX
jqnK0ohWIknhkb17DSRoF5rHkQl45iEepuYww7wR8AadgbMYe+6a0elrbxboNtiA90Nu7FZ2GhSx
McVRSGeuognra8fYgD+JZLhMUqZauPhl9Nf0/AIXBlUvFQg9F4PumQ1FWEmBI7St0hAWlHJUOETS
dHz2NQcKRukolfcAhYu6/MT1VHSMSoJW6Xcqwl7d/jQgf5wWvrKSY4832i/U5uez6imABdSJqd9p
20zjjHNJZT+79MctnRGvYz0m98uWJtpDOdFTkJ2VaROu7xwJ+g96UQxUTEtIvchLaSSiheCCHRzC
jPxu6d+vutPyr0ydgCoKh4IT0CEWEDDSfkvYD3zBttp/y+71rcGnmA4PFeuh/Yc5Y49ZaLxrNW1F
E19wi3oPFGUPE+Py0tdpjfxOLRFfnAHFCNXJiaMaAfBYH53716L4RwZGpipgQfe7cn//DcV2lmyB
N14o7lN0g+Ocu4wJe2meUrSbQWCXkgFFLTwFYo0vEPrnf3KYJ3eEmEPX5DsItxeA6Fbd0DPvtIXW
RH4z9WkcA1t3x6SMEcsZPJ3Nj6+2rrNwpHJdkFAh17DVsVz7LBiFgc+mUi28EE1GN2mDrIXnVfoj
R70QiK9sssUY7cUYZ0/ApF53UndaQFc2eaXvmkiSvVWERuItV3DNfzfqn9Wsz/CH/sxhql357EF/
FmcuDW1MZPIMYKT9E98JjFpnXw6e38vSlkzpyWn9QR7o66Y+P47ogfMXlzNhCTFuwhzWl9xUFPRQ
3Q/ZzUk/jqJHhA3GhwrJPL3nsTipYD028E1oy2N/I+GL55nbJv9S5P1dYJPazmnfWNx9CdCtBPY0
fNqcE5WAjAjSkt9GHJGcPoZTgjruYpwy6Cc1f4Ks+L8oH9TNfk/X64YQNtiWZ2lVcgoRfYC5Pfsm
A+FFeLdBxRkGDaOfWNYawgXuH/2aNyT5hTpsHmwTCcNTyMjdGbF5qjl7T3n6RAVEIezVr953Wq74
uYdGSoTE+yMjw0UYf7+8UthslHgqCb+lPb+4Sm9R7OKTAr9aCgBGoFxTQPP3Az+CyzI/72/uHYRH
InTPE0pZLHFQ4HCo2ATzQEXzSkYQogxLw8Tst+VGoHmQefQCu7MT4tg1gJ99YeDY5T2wR96lDHLq
Nie6cVl5CD8PsxU/J8SrJokpP/YXjx4OlBcZnaxXNJxeraWxQc0v+aXPWhfsG3WQipLd9ErYewna
IguN8fNL8KcdpKqrW+IWGUeulKBJbrTvlOnhYIyANPadatrkpeNYgb1bKMRhm7lPpmPNYtSS7iDv
E0RUpcxDeTSqP5pfseavEKp0xKeNa0518z5p78Pm2KuDwissbYNNJ4l+HWypuq4C/MQJPamJ0wAT
7kBHviRr37uVxYO47v4lhJYizUVzCPXlwZ7DShAqE6r+G72a+dUy7xRc4JFCX/hYDZC9WI6VFvbI
k4Uc1WV9CvM3fD2LzU1bf8u5hoWKm6fCh20FU5N7Gm64jbmxl134xcdj8Brq6HmVJW2j11Yd8NYq
A/gN9nvKYaMfSyAcP14g7uqk1bV/2/YzFBJJciF7Nalu9amQvfqSrpdcq4t3QgXLd0LUrAuQvu1G
Q/9QHYIJZDlA+tCILbeyBx/nkqf58ZlQrkzOiouu91HyjHEMB4Hx0rhzCoJEgWUZ6LrQKWTNkMY9
rFcjBoRnAgQTISRJ6feMDIzJih90Lvf+0d5su6pfPSHMy389GqqqqGTSMqFEbDABCPp/ZaurV0tg
LtpkcMh3OoMfi/6P08i4HgLnUMJP4fyouiLFpTYKRd7DzGkTlEzs5zPLN5Zfyw3GfLThzY55l+wI
aYLufndn/QNECaO7wijXMQUfo/j1COJXMb2uGGkKR+fDbqgkEpsV3Como2QnAl10lM9ymK48PbsS
vYKueIS4eaIq64RDZ2FJmC1Gl1Fdj9Aqg+eCV5e3IFXv6/kOYI+4ugQ6b9pwhkcL+RkVCyOtHZ+N
kFoj13urCoFC5V6mGKcUxc+l6NC67sqKE19Ymmd5yQOYyJC7j7pIYDk0bAthSZ8lCvp/xcAo71+W
dJ733jbZIZgkRU0rItPxtn5XZDwN9VCzLVNBN90z7UGBwivIPGUIP3akpMcIK4lY3t4p50QvyHRp
lGRKRM3Qdk8Cg43aivuB4PqzTPr/Z+S3eyNPo1UhroEDslet42KiKrYuKiLvpzThRuUw1XnS5mlT
4yXEi3lOiXD3jeAUJL2w1B/O4tjBGtNJZBXYlS8j9pukQxTQk23hnOXX571s4fJRyW8VX3FQxkVX
JzycL0jeZQwBCZnpUWbi7isugTB2ZjmL4pTdhHV7cuccVEiEHVuRYVwhpXPcV/tpYoMnj4YUBp9D
O4qiwk61elKjfBS26+zOlNqsa3s3yRpgVNu7BR/OD74aZ/ypU9YdR603QxTfHUyj7z7/efGu6AEC
6GyUaNDSWJhjrDbcgARCkNfpJZlrZjT5SY5t67chUS0yByDbMvwNUreV9dkOMlT6ucKv/6tFVUvU
UXbmlg0nglUOjDdJR51pd3WgJdSAJsIrw8p4+VK8zt1+Ahl/sRWN66AYEv4tntdljpSOiADr7iiK
e+SaH+72xP48LJdnnHiqD4BW0H6qv3/bnIzCmSTfDs7+31o/aV4dglDWX+IWXPD/mt14j8wq763n
A+W16NC9R7B4KObhWtyJ6SkXSLV1d7fBUkLHYY8kE8xrjCgvGEnv6a2I0rWMTym8ielapEL/rTEJ
vO/Ae8/JBv51ZzpkhmmFGCEPUJ7g4DtsymKTqueQxdhlICIvEVTrYNXtf32eoQpLl6kBOR28rp8e
NucwiPfE/oqNSOCOQmkIfodF5RixWm+R7jnP88Vg/VMBlDe4kB1QzYvcegfQp/ATxfaKtD5DaYY2
NZpJ6GIKlRVVfsHZVOw/0/fUz0h0aBAW5DlgOG6gQl7Ncsk/HhzhJHSO8+R6qH3tdZacDqwAazHl
/6HgP8oKNSpXYS3a/BNaIFFEJl//8BSygGS98pVKTxnQ6xboKafbQt2S5pVGgVNUd/vR0xnmrFbk
ttr8ff9f4KEKM9NPmGRKZq2rzOU6+YUh8wM3FHtv1orTSuCFNZOE8PUYu7C/DiHjaHJ04cP2RK+x
AhE9P/h5PMyZtYjjHOsx9nM5u9TG+uteSNVJAwZB9QPiKiff8tMUCKeG7XKx2y6qwsZMSuxtxVoT
R9u9E3FdVIjzTmEdGjvQ1LURIDnnJLE41PT5N+xMHiLQe2dZK4Piejk/3NxrubMuAw0O3n83ueE/
P6ZB3EbXyl55Ej68ZZj+ikLPULb/Iv7W6wQbr2vkENbjwidAPfcNnJv4wKokhcqiGeR6HIVhMCX4
2W1Pd2Jhq4fhtjgTe+YGxt8KPYGJwaLnB784rDn8/Rw+hT5dx9xxr9ggQxi0XdEBtHiFuX7jtoeu
GU0kBeGlK0A3j46RRU0FMDgCurXSTtJ4z+e4w2oE8HYRxpeK2ZdOCoxOsdW/xznqFDh50dmPKPy/
OmoudIIT6LK+R6QEUlZkvbxT7lhiNWwbxWK18NWeNEpgEmb36wD8W/bQ8zPbYvYbWoplpAi+JJKo
WZkB79CyrAmm/bOcqx76Kaa/IC3ajfS8c/Db6yf1vvPjSNruKAprgTf1DH1hSlcAU+TN0BYVIQfL
tjIpoDBZq5C8Ixfybwdrsa9fmwoUZFCMFzHLrARhkoGLDhAb+xY8+NH6q6MlR6vwKtAnsAtyo1iw
1No8cyXd2rn4lW3TV4FOGyTm2DjMuAjPfhLl6efitPPrnQ7kBl23T7qtiaF6CNoIHUZFhmDZhOiq
UVOqqPZvZjdde44l6k45dT5VaZmP/Ci/e2VXq4dU2kxktositVRGA+sLg8CQjkMi3SHDFrHZUGSB
JQpC9DVCmjNRyso3fKdkxhWLAtmqV34UzJvhPMB8Z+t2dB//CSDYS5DcaDMkuo3uVgHSxiXId+Cj
Ti88ghkgqCid9XTl/E7tKlNQPb1ZA1fJMNQZ0QqAGK+TOLgtVKw4eB4cbWaUWITs8+9PD0Uu2wGD
eVRXJ+zZhk+IG9cYOdnZEEIsmocbGSs+E8DhoBk5AicjWlfPkQqOsQyYHElJqMjr1V+AY2Wt+FIc
dJAyRO+d/Z9IcResK5OchL+ZAiEew8vg+G9gtIElRMZebIJXoyRbov6qPeFqAsS3VKFJQNJKbQci
k+jOS+pNETMdGFfbzwJzIrX79jMo9uReBNAn0w3fs3wwZ0GvSRELLGo0yPB98T+zzM4ew9cb2aYP
0+6vrowKmzNj7AE8B4nY92MUUBO6ttWy04f7mQ4cdj2vSQ2INeL71ZTFUreSfyIY9a4UXZpJK3Gy
s6rHk6clhNWTnwvRScIVgmP0ufNgpXFBS/f8wnp4tOBDQAYTwHNSlf0OBukiWj9PyrrViwVfKrT2
2fUDcyDudjX71ZikFCTHz2wGN3Peo5mUp1h/iC9wwEF6492ph3YbGe2z/rBAXoEMOSk5kvhVJJCk
WXxD8yukMA0tV9rqxrJOZCVlMCEmGfxbOI0tIMfsfS1yXxxrQ2Fip6A5ia2TLy7hnlnNF20vyFJ8
fpzhRnfGQ8qkfupGqCvH+S1AfUw0k9WJHVWL+8qReWORl6G5ha5IwA7LyNVD/44lum48jbFGii1h
aAJSiwwnDr22QLTWs7SmLCxLqh/Ttpwjy7s3gdaZIVUDxUQzghuXyZOuXza/L2hRpOomw4JY2fEC
ud37tJWgEzsA7ubdk79OWkTXzdDrMlWUAb5FnBhHVYnmZBCNY2SkVOv20ZsLDm7dl+6cjS6atoFJ
tdvrxlayxkK7gLWomg8whxO6t4onfG1oi3WdQZAvRnoVUuNOSXZYJXNLOD3UFYd3M3Y7480FY0f8
ZCFrWUOp2o3gHb0vrMD4JzjBTdCMqIB0N1DVDtyA05PtO5vwj2rWLYFtGgWXAKJtoz6A/Xbhgp0F
5RQiwZOJPg7J0rh61qBg1iT1QDy348d1aPI9Axqc53MChZdGveQN2LoDCzBO702k5mQVrp8ugZ3f
2jT1LgbI/mOmsTES+hL7PfI1qJt2xILkOEOost/6aA/sgeJ3SqF0+LzYusKYGGGP4BHDQLRnJYuP
wgCI4wuUUu5STqpJxOMDWWlkKBwCha+0W0C8JXiayHChuqFKCg+mt7b4xHOFs4Cgjn2IGbK2xO1F
5YqqA8wxePPT/gtLJuKyAYYdeHtLduAo/A8Tv9N6V7kkgH59lABTQ/7WYKbmw1l8MBzy2rpko9g6
BbhsmBzP6oEPgqHV/X007i5jSNszWX8toEAALvIjunqOwWI/ZgWWZLO/Dsnt+R+zQU/O9h1JgyNe
FuxZw+DyUH2OU2E9AvegCyA0+6bDCkFgLO0S93Y/pukULTts6sGehkDzk+6DMsr+n6WXW6iqrfw5
n0xix14Qwlqf5QOrBfijaVlJqmU3nPR7wq33bNg7/bqCZ+JlCnxJ3FFXx0Y+7JsyBdH9cknwEiMd
0QYBS6YjV1KDXjs6TKmYwpVgzvZyLbNYTvLRa47+R0+SmJ3RbKGnwDTAKfwqiDqOctPzXuja/zCk
DXkqu7OOoPcSsJa9fz/xTFtLwANnvXDw8kY+rD3oTMOTTIG2977ZcKMwW4njhcjtfcoI751qXI3z
vuawdvkQfros67clT0myPylZTPxtm/9ECwrZmfwYoRkGPUZjE7wLtThb/ZgXgY0QqL7RjBq4NEuf
PLdJSBNII718omHNLVqUhh21ZCgRWYgPy3ccoq0xmb2U8QlxrURJf+fu0jirNlHGpM6z7ma5IIH4
ZBmpa4dh7DgsGfEyInz+C7Axd4NrCHgo9wQJO3zCeXIgrUljrz1QG8FeZDkpHsRCwxT1opNZgAGu
SlRAeg4rrwczdOSdYdr32VVCtfL9UolLCWKQZj5Ta+23IgdSzCeoUeubLVkB2D51Je7WrFJ5rwcm
weD8a06DBDee1nETk0/NdRBVAmOo9wSs7vWgziEa307Xbq0RQ6mDDj+WqA0KRZl4q7h0qmHv8noE
w5j5u2Zp67tRQCnkDDBpUlyW17LrVUIo5ZrCWZQed9HqdfxRMelE3d333zUXAIuYbksynk8DlQJQ
STfWt1wy54vtg0capKNnexJBXXJGgWqUtLC16MqvuuUGiR3DTvjka8A6jWyr2LfVQk5w5B13+ptr
5JGckmPm3HYre87lfspriSzXWVk5XPDw73QpUFDIP/UZSitusvMbmYgj7i9dc4F0HPmixVvvTsNc
MPrKAkr5UrXfBFttrkQ89mPRpX+gtkQPXfQdMOw3RUBNNK+XasngTrAEEH7EgNyPRCtiM9GAVczP
i52njSTqOT/OQHn6gICC/44ekoIsdBMsZGCt0BDmws2awyrLW2UIDd0NsysIy3lW8osh+28pbvW9
Caw66cNmUeaK3LJhBM1kimEfkrerPmiXmFJANrfT4GYk7JYB5iz4323pZMjab+I81zWMyHn4pFp8
/gJiklzhunAZe+t1yhzXDOojuzyjd20gS5XL8AODE0Cxeq4+/7H4pdcF+cdn0wd1jUTBT+12kInn
WDiYQk6VihCPV9d0+6fA7s1UmIJnylQeU+SiIwfiCgXdm/A9tQ8CV7ot05puUjS75/YAbU9V9xRa
iBBICRaHUv02bLj5IV6h4Cuzjd1s+Kj2iXSn/IIWAGbYAAUA0vEM7wSa/pYrHJSh5tZha+9Q8nA2
ZN6oS/gOeqoyDgaMDCxxakfQHsbgLs51nRp0+D9WlTG50twMD2t+t4pxtQPhpRzw4T9NHHXnY437
270KakoVpZqzZaUctE4KK5rcB70JCDJEnhGNJkjIvcTsp75+YtY58iZk/84bV7p85RPCbTHRTPvp
tN7xfPyXhj0twBknJ3ti3Mm8Vklvp0/sFiRUQPMkf726BGLy7DSvdpuGX/J6KD+1ZzUozCKdW9eq
AEgzG4BktqWTQ+1jnoGB3wNOsON4Sw0XNzYbWEPq259GoKtoOKv8ZoLzYv0A7qLFj7T/0Z6nI1tG
7Axoy0maJBWlRY89K22rrSrt2VhGLJg4SuLopv2f2RZgJkaCDxAGzo7ogZv8VTs74T1Oo3P8Vrx0
VGls62PucN4/XKldeer5ND4gl6jed/S0WKV6XGT7uvsPoh+OkJMvcrbTXREyEvilSeFzs6mL6DFb
7pliqfU8ZhcLXsQeFwwP6aHxFsaKD6n4uKgNNQ4OoFjk1fYCULou0xzUJdqdavp14f/XMb8tqNmM
+oOyahaLxKHXwsnn5CsiKiT7iSxsOIace6N//gfkFdna4wcFutEsByZvTIwWxbhWszxBbC2/Xd4F
Mt4bIGDgoitl10tlmIHC1+91uDj3lKxZXWpDKl7KdNfeNhP2rEfU2YQuZGHJHPG6hhh55b9HLU7L
Dy+efa7OvgzHbOR8k+gPpw70AJWc9uwy7t7oo7QXz8bZvU7fKaCwl6niNdJo4MVTiwbYZYOhDowO
+unY34oqnE7Q268ubQJSIRRUe/DhXlspp6YOolEXeMnkHL/Uo+joDCbXazyI0OjsEMWTFtRocti8
Pwcv0amUtFpbVSQYdlPXlaYlpmaC1nPtj38Cb2QMyzabis4NsShQZouyfXf96ZTgCqGP9hf1snBB
X9sqrYhcrU4cWgRiuBVSR6+WAJ55Ri1ySDw2oAhVmufcpJbOpbZ/SENMh3+Wvfrnr0bl+gj/xij6
GnQR0/zh43B9ssalcHuSm8zh8nRQQYfhCULQa+mqTGBwD5R7aVgGg5QjTw6rpZPxEJ+POwLu6l+a
6YcZqoXu/OIrjZbdS9Ny5nhwy/E7uXBZ/llbWNJeNc9CqoxhIGiQ9OutTjESU0AHpcJTGhaym/me
gGS10ko99AwaNCElGH2bN/xs5lya4HEXX7OuVvuSYEGdXvT1/RGYFxDdOPcysMCmK/AtKBrataJU
idrIYsADZWS2w1pUJhihTwjEc/wsvhI4DJ+fGPg6GskYqEIaxNpvU+dGUAHAy0C5PaSdXkNzFxmo
yjVVxqx4SwpV2pvYk++xGNo94km8d3nKKyx8d5HBhvRZ72sA6hLPUi3Ewe5XRDNyobJw6dyC+acR
mWOhS7Q4W5eXfo3yOzcE/gMP75QLVzOteohcXFBCavpwmIQLFu/5lJjJqoBNxpUdaw18HVjzC6PO
hZB4MWIpem2I1NY6QLFLR3hj/5xLaSRhRBsHuCAqFZUDhXVUOEn+rIGWxBigI4qoTm0MxoBobcWU
geupvNHmGCMOl8k2oMCieY1yXqEltjhtwIoIG8NQlBilviUaWVk2JkBcsFr7HVaeZCx47j9bHvAI
q/nLm60O/vlz3OQPU8sG+GOkCQWJfhiQ30xPuKbGlat3bCmP/ZpPrlbT7T0iE272gLc3eE+FhfIB
KOPpEmTnZh2H8ArvBrxD7xb8aLRV+MMWSDbR3BaxluSQxNjwzrheqwvs7CCiwawwuktavvkBqDJt
C1L3fFHQ2HV3QgIR/YTY2PNcu/FzG7zz3h3W6fJUaN628p7Mf5zsWDqoHw4rKZmXhISKcmsjm8Jo
1l3NJubC/+GdBsK7Ksht3PlM8QhGWmq+ywBQBzlTpLG+lg0Wo0DyTMTiOzX+h227aNuJLkTFFvIE
8jr3LYhygRqtkBi/92CKqS5p3Ls4/cY353jfENQmKilU4j/pY5bwKAxsbr2yAKRWNB9y4ZC6D6hK
O5WJA1hwoqQ542U1VR39oQojGU16/nFyYsQfHyFiZaizDVM8KQ1Q+4Jg9mJ4DfeFCSVmJA7BbKZI
57SDVL/oiUHJjpvqGvlTqLdjzrh370y5dvw93hqBcZXsZFNCbS8ZxKovCySOImGiT5I7XzwlxC6i
GlVDMQrYR13APXHcZfgyrMcfFbuykjMseVEXGIjLGi9dNPV21NCq2OgPf56tQmCurxDP581VqPa1
/quxKp5DH0t9OgrvmFZcaUDnvSIzXb9YeFe4jSK3ImQhNTxNtPfijalzXtbMIFo/9xLa6qcOyZRw
eux+AUV0KRTwQCSd9GFzx3PHpLgep4dTU0jEIA48fw+MElrKZapgU+W8sctIjQA0PTIoy/xy4LYj
+xrr6+BLWmXy2stCDLGFFG6hzSkHBxTOVS8KBFRsYu0VaQZ2qyeqUMrHKCnIt5LFWl9vCkwcbc2f
5XKPL2/jh2eog2/3utqDlDk9xTzP6O3idyLMTeRNEv88ZWeRuIVceGhn5FJmSp7XoPs+VuWXNEhU
on3I4YGw9kEOKHrAHRcqqoOp7WcGVZ6oVhkeKdekgF/a+wbMg5OJMJePFLe2bg0uXLgCObNQ53Fu
c2vaN2MWf5oYDoRZE9dpwW0e7Ircleb1bQVWEypQY0RAEdFCvRxPhBqRBD9CejIuSz3U/oM6RMMr
U4PYuIwZBk61YPnt+4CX8HUj+RmXa9eYueyeKqax8SGOO+48yY8zwQPs2S7/zBHJimBLKOK3of3F
t3Hz4OVb7RcwVroWHFTXZVebzZvCSO9rWFOtYbNgdSpAWaI+Z6v2yEY4mMjGROVcYG7ANt8DO1rG
OJgw7BZ1QcpzeRhhDFbvUW5IZ0EEUgjduNfxoggtYixJUqdJo0SIzpsb9jg3V1WI5Ar6Fv9XC+/4
PLUU5ipek9ZNRN5H6ywOmhKzeW9xQRy/Ms7jrdfQiLj/dkV6HS9QDZYc+ghkfrrrtoiTNIfTZYnK
XL76nvwQAAbbPW0TAMfhYhmhEAjIoS1Al3RKfmXOWIEKnmGzrqG4NHogWTnpWeZA9Fl2Xz37qjH3
Rb3gGvdv7IHob88LtigIOiaA3ircmIbb9RmfmXfcHlLv6hABjneLjmBOQiKIMRGZ4yv2YfdUCNBi
D0DyL+E6a3I2vZj3lPJ0nShJDLq5WtXBBUkjeouMpLSWoslAoojJMXtmIAkx7wTgfj9WjuLO2zcs
W2BIJq3omGO8In0laz4rZXSP22n2eFuKB+Uk8kOdfid/zu6XjQdv0dRIhpTgEIMUuGWobNNjH5cM
wtwWsjlYhIn3pIOEoc5oVra15DdTkpSR8k89u155YWtz+IQIw15/k3uRTewljxBKKd1FFITGcD0P
JfB8DyYcfpwNPBoAlGvvI528qyfvlKNPfne4mjtiz6tGwTFkjqaylWGWO7B+YIEEobKGLePwXLv4
0RVxdp+tBxa6+mLeLcUOtBumsda3siMb/bHrU3hoiqRwtMw0EHSS2nX/Veqy1GWTpRmhHoMUDVKR
aDqyNGXpIbbxXsGfNeYSoe5jZnD1O7e5Fl6+l1q6x01DuLt/COBtTcN+D+kb7doxkb2Wq8AauarN
Oalgu09rhE2c3V9R8SUd+QsJAMvYTrsa/Br2tNawDyuUQ8+qAiYTXNCrnxz72/bWYpoGuzy0yYXW
Bp3TBTs70wzGChHYoOCM6cGTEVVbWcBFQCMzB8VfKiQ98YqXsqeRA2clk58VmqJ/zIrEaTOgviDB
CKOruPVAvUmmm2Uk61Zfwf46eNZrNkIrWGXByek+Q5o0aU9CFAQcmRp7xxn/h8OlnM7+VATugSx8
p3s9WIste1SqAOydB9lWYL/dBXWUNvrv2G9zUSAJvyO4ygznK8s+wjr/BXo9ibqHTm8Cp8ohXsf1
Ve7Gsmn5fU73aNzac5UCguYTAQX1r+2mjY0XKTwN8h/Mze1mKqsTj5v8Xu7c3zu7xeENkfex7lqo
W1k3YPt0gintu5Vlgt4mNSXx3dOd9PXzgpNiSDDfZudOMFoEVqTb6ppKTay8tBcSMjtVt6EftbOL
rfUV+d/zNhwEIQRbCpRAOPr4HSA0hL8mBWsDGJ937QLYf/ttafMlKcCZHZbYmhT5tBmCXtEeNY/K
r+A49phlM6CB5NBQZ4Arugdw1DLXslNBg46lrfuWYFqCjBiXznVA+LyM5No007Ur9Bqk39IjqB6N
c/nKmeLslLOGtuat9drBL0zSFZIYt0EPSke9Yf8gVcYMLz2f5MqoMlU5G9M66G98tR1bF8icIuqi
JGZrmnaRcIEQAK0ug7B8bjMUT0c9SlG0vRsKrjvW9vLF7LdH+uPa+OzQmWsxyfmEnROAaNZPcwPe
UrX1yH77zm4AlBvAYlPEvqh06tMEpmI+DPTkPsr1nu8Q76RSTJy6y2D5SaY5jtNLSlv0csINNx0T
9UHFhRL0WoVdYjNC+bulXC27AO1FqWV3zBMrMyWV3sGE3y0jotohvhIVK8ple4oHki3IiZOlMFvY
FOHOThfHTWxTKVZkj7UWs0+/WRNIc8dxmPBsCSg3mT1fGpR6BIq8vS4jVBN0hQTxMoAED7j5Ie3j
v+JX/rKXmcDZu1bRmiUbt4gsElnd1XE6UT6HkW9dsLHqegiMABdawD95egTvohUokpRkdaD2GfA1
eEH1C3ebxYBmEB5mV09QgjeCd4V0BS5L5TSnIWpZkJNbr2XPBoSrM4Gagdk/QmWq73JvyMzEe4t1
itktt1sM9zsFWlYVYyh7i2zA6SZ+8S302i9WjBbRmdT0Dy83z4FeP+F1MxuuiqaiwlubtmNopjJT
wtlMxSoNI4AX6LuItT+M1+TKv4410gahrzecnY+Uo2Id0D9cksppLv4nXfLA1oTteEcgswLHsOjL
eHPYsT5ItLoLS8zm3z/hQohRQRumgFCsDF0kRHNPfRUdZJInyaztq3rdjWXYghUF9uhE9SIVpAME
VsSAO29+W2/CygwxILFhdiux1flseAZW+iyBTZJkuu40cWAkfb0dgS7dOeEu5RFQlp3zshfXzmEM
xxx1D7z3vF4TmkxHXG5H9W3TnudkqBGrJ4ijpFrWhjDnLUtMLdn0OEv/wNpEe92eedtu8wQ5L2of
9Qhxu/mogf8MgArwmC1wZODS7KJhlKnmxTtFREKmIU7JMwNtIYKYG2KukUMWyhjVhhD0tMm/Mss+
k8qdqIOV7Ey1+qZ8aUCuHgvYfnal74uW/mtVU54U+NlAIFmpXrLVHzpyiIWAySBeyM7PizpblbBb
53dRdAH6JzeXl0ztb+mK2fSk86WNC+G68FLM7SscKu6INWIvcdAuY7DSAfrKNvd6sSYx4UBfchO0
nTtRyAxjSzCOsgjnTgPCoJ6wrY2CnYrrx5tisT+isjMWwvMR9Z/WVHXXbdW+WuC+VcvpldjTJFjo
Q/cZPScJikoqT7vx5F1uC6IKREiRI4pWps/oSuhO3Q3c7JWGSKKLw2lRUxCrhBdBUEq/mnhGp0rn
zpcyRj2BjIRD2O/v92aR8vA+E13mlt/SOYRkfU0Ok3u1/IT3VOqdklrapGcvTgGqNtAySzehKZJY
h2wpb4BamVdDXHFTXw/8RJ9TWdv9sJzeKgCyTHYdzXYfNxxjb/WK+Jwo/Rd1OJay0XLzLGJHG/Lc
ks2L28N936fj4uyJ0CAShPgNEEOjyOjqqNeMyHlORUfa5iI1wZfxS+saOw6OXtCGBxZtDEd+Tnes
eprtjKG5QlrS49a46o7X5PlyXmIWv6DaifM6d4clDq9wk60jxy4cJLtcIEU8666G5Mdy9TVOcp9N
xhmf+0+sPm6pGoahaUfEw5wNwW/0v8+oQaabzRY3wcfytX+9Ukdj0/R3UviWHmQ4llgqVvAVMA9Y
GoKH7R/suUmgLA60XRr0JI/XkeGke7N4XqrSj8CbWdXOIzTGECHfWCffNdNVE9MHOaIT5BqpW1Pi
/+4b4yboRraaSzhZbpZDZ4Q8DliruWSnB2/XN0d2wLF5EAFqw5hu0t2p3dAcBqqklCE6kuO9xP5y
7COuKuYcYM2StZ8tLl5DBGGNjcISpuKZ28s/7xYbplHY2J+AN2Fw7EI3GKaLwFu0HjlVp7IrqT3i
sU7hTCXQrs2uU7nZqKce7aqDXS2eZBlGvwVBhKXcX+37o7WEwj70znCWl+SpoJP8z9LYaAfqarP1
cPasEPAgPa98GjgquhHVO5W+6khM5ZiswwFNYC8Dr/D5HgGh9cfEGvkG2vQz+c7FSWDSVpxUO5mN
9YO8uR2adAcnMWWefq1QGdf/f5ZVpMrt/NgSXcaYcbi7dcVa3dQrzaA/OUY+7tVq8uBfPXqJp0Mb
9GWLzaVY3tu7Dq1Y5G7McvHufGecxa8KzDEyKbKSP5K6NR7/qjj6cOCHNYuzJJbn12xza3vdiuks
DnJ8BeQRgShpW7jOUCfDpOr7SxyayjoWl7BDcQtBEObSytH6qH/JxDSisX/I7LErIHN6uYTdFkBB
J9/IJQ4s8fGFhkQMr9zFrtJ9sxDhUSUlJA6Lq8VpD4hxBIMZ2klriJ9up890KHVx3D1deljqvtZM
84bcXFMPhn304S51kPor9HIsqxqUB0Mjoxmgbd2eXj61RKhSlG42Gx7rlhidJo2yNoEESEAoBP9o
NmDnKm93zWA1Z9VhBPRFSs3A/WA2MymImKYfkuKdKFZupw1xdEbnfOZeMRUO/ucg1za4H76yyWz/
DGaZ2LzIk75OPoIvkrWEQ0q/iiNUpEOesgaNCb0NowD28nKv/ajRRtf4BwpVs8+zESVuHImUaCL+
I5DyVKBWY0DZeadsoOuXdE3/3DRaNG+kYg5nuf6y4B5zrhsYcXuM2rsksKwHB7WElWjO4fTu21nk
pxFuyLIdHp0PxrlM7jrBLkwcBKWJ27DKtBsPT0fW+aRHOxhJQ9RxbTxQ9ewRdxLbIS+dslG8CMkd
6wIKo0gJNqhAnKtfes0Zu7A8ycGSHFF6TphABzHFa5uJGw/gHdlDRxli1z1N6HA3VBGOPuJmYt7o
gCsOPnClR6lipDW2mxU1Dzs7Cg5kK7NxF8RdmBS4Q0h7lUMrB7cFr6DHtw5IfxUWvap2rvSsOUbB
+E02mKQeysZlr9p3qdTmVAK5dwtvg1XkUb6e9gL+1ZcawOX+6CF+rj9b733dlTMnUae27MK0s7Dz
9QlUFHv8qbN7GDiV6SvYR7PPEc17AOqz5sKNTeGCOwy/Hbx/eN7qv0MKm5X/lNfYB4KKYKasqacd
ucK4zW1lwFOI0HT3pZtGBOQqlb4lRz54+b/jnuaOwEGRgH3W3XuUT4OkZtSf0pEogEP2mBdZrx1J
JrpZ9as8xCiI21mr76EUvPX/Ch0DXd4ZG/d0MxHEYg+2vD0esodQTmRnDXHl9m1V80CX+vSsSlWM
V0rxgUBmJyOcPAtvpiCoDYu39eVBlQuLnJINYziIHalH5BcdaECvA97CWpRwB8ZVYuxymWsJSozx
nKR8+vjvDXUYlrKHEMsNSDNdja9BADmFExw8XIYmJfxVUDymw7KJ9CcaNs/kqqehATUrUot8Y3Me
d4PEkZOHKPG2M96CN97ByA1fIBn3HV7OixNZ5Is8HajMHLjz9oQpKrAmqXzwoph82W/BDfzkWDvX
IdmGUe3t/mpg10CG8LvnDJXS50uEgdbepK3qQcyvF9h8LislapAHEV44f60XdKVi+8LUYx8gXsvb
G9YbHirojHkXsLu86iMlVqpsmnFM+GqKDMwsaSm2u6GsqxedRd9j6008KzCOh8I28+3jq998Pb6U
tJoKI7jfaDqgQIWC+Fat4W23CkUac+haiOqN8UCeY/36C+Gz1tGXJFtDfkZFN8Ui41SfHOG+vrND
ni+JsstF2UsvndUuU+x9oNc6+Gqb7qICiyKzXm3YKJqo2h2jJUHk7ALMCrmio/I4bbi6kq+7me4H
4Kbpx+CQaV2PuU3hduufBBZgrKXPtKmtYLX/DkFZX8CeOkl2KZ3ArVz97uRknXa3m0rS/QpaV+fx
YPIAamZXnmQU3tRfZhHmEZRj0NfuLypvdG/zv6dS8ySDYnA/pV48Hyt05PdU/svAmOY1p3DwnvbI
4KXwVHt3OpSXSLfr+z95D6ORLfCowQyLoAOb7rYZuKmv9v7dTUwc4cUDufBIltJ6HOc6FNMHYvwt
GBA7LNAZVw7LIjeYQEBs7CB8zf+ckkNxnnSKfHoBc35jT37yMpeOdjejysC6jrjY2azVyH/t5eKz
KJbKAOnIf5jZezRUhpeRQzOiRSHPsHa4ba6gjkU0p0CHsd5aTfLyq4l/ffB/3/9tD+4a2mVb09Ft
GpcdBv4/IeJ2+DsmRS9pPSOxc94xA06Rf+aU8UCfCvAf/yeM3ZNW18qucKPwuU2rFnemenGQhVxp
h/5QnAi0jVyFMgI8Vj6/pjeYQZJeLD+05P0WLlaaAfq6y6bFkClA8n7GJpnLsUaE3UW35lVMqUEk
6sbvRGjcdsYjb+y7AsNFHvHLA2z0hVQ3J5WfTboDmLy+Xa2F/0syYCjMyHxF0Q0nVWjI1CiQpzv3
43LSUYBF+fewrqSrt8dIPD40W79+DQOLbN9PZXwKIX6kEAvOMPtKae0uQ80AvF49dqWg2kQooRUE
wFDTlA4oYMyRyDtlhNSE0+VgiOLFb1IGS7llryIfC/30LGMH85Ju5Vn3c5cV+BlCSNUHZtHuL4sS
yYqXxyfHo5+Ja8yOXpVymlma8bj7EOCbrKXoyabYXoAcsPhQIHQuVKzIrul0m5olLNM3TqlEzmQE
ykLy53rXxQNkUcNc9Y0uUmKLTESapxa829VmFT75GnPg/HqJwFj3q5hPUWvbyPOyH9/ERqd4IeYc
vahUgWzeLrknoYakVwQq7KVf7X0rPPvjIvYqVzqo6BiefZUNzoUM/MTiSL0Lh0o+E2ZK/8hTEgrL
nPMPSEXw16f5KDczse8uGX/L8Zju47sD6Q20WO1F5spwWmoPLg5YDjzkltZ64XI3QKJXk+Qk+f6J
gB0QBMhaSqV7vEecbrU4Zqzvok9D0YM60KKeaLmVRpG7Es9htr/zn3ofsbbmXuYp/06KQAhizrnh
e1MaXvv7P5Ucr32cdFLhfnAdOinNztXLFq4ECL9uYNngWAW6Hpx57UtKYglR+GciaVge36d+KKMY
OuEYb9MGWs7nOvFgqu4VcqiTBmVQb093DRUjVWkbSZ822wuarCNJqv4K/xcIh3hOWAmoGp2+/Eww
YQCYDj+AIOWSa9PQC2EoqO8SXv6VAsJjqKlgVbCwDamHhYpnGwmUAJhrjgRgYxBmzHaiWSA+Krtu
7NLw0D33uiVp+ZNj27Q16WlJWsxENBnhgaoH9zdEYekTZE0hztOqrGiYcerDaGkRQEYE/nLqJusw
K6pNwg+i7qLV649LoWRmlBsJTLa8IoINxPLxQpy0GGk/VpMDntI6rfj/khD1NefDgRRxpXNzBzBI
DsYNr+IOE69PJv8z9exvQ+l7Evmy+EqIQHzGFNtEx1j87o9V9MiaLZ4izZv0+C7CBoQ1KIc62HKo
T7PE+tzQLQBQ85fDqNRbeJ1Gp80CedP+heAwfVxo/Nx1DRxjcMtA5/CKr7KE4+EhKYFvw7yb3Q35
dFGdIdLAnjpGEdZdNIBaLgLfq/k/dH8an3Afo6G6c62X7nQt7KDeThOkAbWYSyOqRqwFtpJSgi7E
KzeYsiJiNZC076Pc6hVI6GnyPAPe0EcRi+IQfS+eo3GhKFjC6EmQQwEW4nd4GYtbIrfrJDBhlQXG
1ua5t7WzgjYCmf0oj5qeMNFUP8gklBGLLOotY6CdpJCtdjxGFv6O5EWO8vhn6JdGYk8vRDDtDB0L
WGQEvRC/AvXqYK1y6UCrVZ8B7oflS/DupgZe0JAUPEtLhQj94r0ov9qgqzPhnVMpNSBIk/nlPMfG
5imK1fq7ATbJECl5E7K2qua9vriCjt+1n+wPHGRbVDUwtoXnInuO+e7ZlcpQ1yg/H43wZa5DjfG/
YHM/SQ932lcLLuIGC3wJkknwtUBdo8nE5P3HQPhDAQlONPqlFDlTBE/cpxWSbaM5+ypRB4gN8mRW
I+3Gxe2T14oLk09CIIW6rdClxCMD9B3HNtzCjgSLDMVmPn4Wq1gMsxyXIqO+ys4H5tKF2iY3pMmY
e3hCJI7RbA14nevkJWUui0Rm0VWS1yK1JycAnRpkjKc9YVeA0IvPFJNzXs475i9zqRHhbjVQ5E3O
e8KWxswo8Bj9M65B6+OT/aBUhGvdfoKE7cPnq+mqMkyIbcCJiqkG5X79UJ+cBb5kT0TbU9h1dEQt
cG/L8P6xDYMn6gh7HnnLs2VlAI+UptVbqTp3BZKlfRbSyoFn/3cX2k87QieWq1l53EoTNKxTA1Gp
Pdk95I0Hl1igIC+FYC/SjhII0cNFbuW8fP/oLehPp8QQ/Jdc/Ypgxf4e9xB75i7Czewifqo6r3sy
2Z15tjtzTvh1/ZlH6rVm9Z5iorYrtEJBb3yhsDPxobPguIEaOWqkCMV3rUG+hrdi3dGSQGUqlCVi
DScJ4dZs/pLTP57SvoZ4CU9eFKkRMcILL5+L+q1vfHWiYVR8ND/8gHDLtjDzA/0F+VSavUS9WFNy
TVmurOSaH2rJMaZBHYwpjj1drlC3GNNIYdPHoYy9abPxxwU56acQAssFo1FDg4LKYwl2kOBu17Ar
ucdpATEePn+RYxIfmfdAMgHN7sk21shawp5rmGXKM6jAalj4uYZ4gSq2+dYV8DueHAQnXV5wUnro
lPIbyYCoHxjedV/E7wC3W5Iqz4+DoSNZEPDYWotlLuwRT451B2Hkv69Rufz2cDW8j9O5VJO5ksCu
BjzaCJax7icE90gs64+sjMtirDe7NsRZynbWY4aN6+6RS7AwSRTxjPXir/iUDu8z7ybWqNeq0/tk
kG9dtikR7j5XkK9a/VMdCd/SB86ySssLDbO1KzC+h0j4Hkm41rnxRAgq+ZDIQv6nbyoj26cVnz/j
Qh7jGJ6k2iCdexkHHg4cNPUssuMRmP752BxF90s4UTUsxgc44FNXqWGDObkaIPIHgw5KnEeLQtUO
MOBDx3BW4doM5Dao1xCRqHxM4Atonj0Y7qArjjcyWajao+dsSoQhwBrk3KuGeEDNple3Vco3hFmF
JWCmTGLOArNjTs6Scl+z8pBYPAU1WPxv7eaeKcFuR2lsTeV/kGjXif9MFv6u53Olvtm6uDt8RSa1
x6SulhsjViBJSHz6NiIuK1GCEtbn4n5Cf4eUKReNOWrwEaKMgiPjepVgtkDnvbM/wVhj81Pw0S3+
tD1R94Y7oQ5AKc3AJYwzbdhDXM0wakpJ9oonue3gxuNSXCsZvX6snvw59qyIjC2/f6n3OlBkno0M
/QrIMz1bjg085kM7FRpduOQufB8xBHAigLVIHxR+G8kRckmZckjAfszk4poU24MiazBl4tMZlpLC
XCvkb/5Za9j6tTKLRBswKF6LwxobTmteYdEDEy+L/n6Lt1rpjf1KOQ3xKrsfJlawNFSR5d69paPR
GvgLJkHf4tqmw8sGObabbZ8OcLvvfk35m+8BkJtrOsIc+4nKbY2UwODyjBRW8w7v+/awCbfpxFL2
VZ+suLDqdyGW7T2BR+KTRuZJr+4VHAp0i5ztwKLTfB2OLbP0TpANo4/ieth59GYRoRrscj3f5GtD
wcVXCwBxdpZ1tot+7A4KlSzUqA+xtvdKSN5ZKgk+iuQGJMe9xtSdCKyGl1oxEJy6HHpJ59jRRwuq
5IkN8a/VGqwFnIN45+4XtlmmDzUTmwrfFD77cfcmep4iVwWDUpXCz/c/pDKckTTNTVE/j5bIhz3m
WYdRFopclMZ6wBIkOToCUL/YV3tzQ/MoszINTG79Qq8wujU0I/xWSzMI+2ss0O4fDw5rP2R08POh
0W9lF5Aeb++ZpYbFrsr15cVMsLxmlTBouuovsMQh/66znCnFVtuGT+WEEY37LJKn1HCRl5CEBtw5
TOGLXcY5sxMdDcv6CX6LSMbhDa877ZhM3pkfgNhWyzwX5mE6mgZej7mJRl6pGOd1Kvx1jCNyrIro
RW5wJXejwe3Ri0rhmUFCr468rF73y21a6dYv6kPlxW4pr2LTKvpuf6bCqLN+FBus6uw8eE5zt6Y9
Ww8L48bGQcn0kpWrxl5GV4ETIuyMZ9Pk3wAHH1tEJchZt1Ynj3rp3tEYZxZ2p3R2UGIa1JbTFZ8Q
qk0pKUJLvPjaR5wAZKVIOX4Jc+W1O8aobwcmlorBcVmBW6zr7b86m+t1eAAmnInDHS6PTypOogyB
s3dbWveUfXMHFIExmi5hyhlp/fl5e5jdxRU72aDfOODKCqawYyJmppKVNW0BwEuDQ0F36ZygA8On
SeP03s7o8OqNTs+dDHPiXFTaZTygVdf07Y5u5swX0uIsaYqSQc68Jfo/xFRDlwy+zjhVdOc+IWSE
49vIaosMe3AM42vP5BddnnpYB87hD8pVl+fc2lyePSegDGaHS/SzzUQXVKgox78weBWKcCa3u3Uz
F3I1ums0XO35qtZYumxuFvede7nhx5dkkDqXxNKGhoZU0yxCi2SLrjVjlvtw58iExV0gxn+/q9HY
hN8g5085N9i9x8zFA1PZwEZ0mvWXbzmX+JKc5uLGHC4xW9AWLg0C90oRZFXceRsCg88wRMBgT4l0
T6O4DTSoNOI88QeHdG6wv6uk6PwIoOXuFPeiJgTOJ7xQ3asRU1qinVeuvSYA/89AeblbyekUOfui
4dvlCEYTeVuBYuAgu409mxr44D7y4r1y6iXdqvxrfbE8VCpe42U7xM5CwQ2vfVsaBIVLq5l4mV2O
P7G4StMp2ivCVpYCUEHiBchy8nwY67v6yhXtqsFrgipw2vqlFMIo4D8ZyqTHOzA3LSEjp1RhfXTO
DKMO6y/7pIlBDIFKjXKgokupjp5PQ81iA6pRdCTZqEFFSm8C2d0Rl1H/OrX+lSRNYieAlzCHW2/P
fbCwdpTz+5ocB47+6XzHnL5q9qrqZkcVK6t6NpHkRFyIRRPBRIny9h9WCKywfy/GYe2P3zJQGwRY
cn3h3rVEe5lmoDa5IS5KWBUCZRFgdtsbIAK2AK2TS/Ng0CMOIyr3Qha3+mfIpaO8alssu0c5g1Id
WEdpdnN44G6E4IggV35hNDvLfQYINupAA34yQrmYCcr+La23j+45kCmLvFKnA7BrVsjL4WEdQG63
ci5HmDv3FFPTiruebzx5gxfwmS0aNSLEa8d4pUHfPGibN0p+K4MG8V2E2m92ZlgJd3ylIbw8QIQt
jxonsIrK2sxkdHuILnHXvMD6MQ5XYwgtHgzuFjWp/L3Exf/WTO84PXq5FgM/aEMYymua2veUy14C
/N5ywUB0cLJdh4qmRGAaR1BV00co3FgCVizvX9tyE0boCxFl4cblPq1JPHiC8lxngdeQnvi+9l+v
7sRN5moa6XHYAIxQc21G8pYnjgK56ZoDPXpWLiey1eEFejvVQJDqpQpsom7sws63WTtU4vu+4M6R
VzhVM+ehY86M9fxky2AWnoRm+N+DS6JXIad3ovfHRSKRMAiaA1KbvFCXvjWPe4MMh7yykCsCLS8v
c+55yXFVU6n2L94bOJEesW87KRjt/htuoxLFk2CXzssjEsXuifCuYOss6IA6cUlrUrLt/X2895aY
CWw+gpkYnLCtiujXsmXrbJj6Mjp+DGSUUVe8FW6nPlMqewehLGMf1KgO1Yvh9nfz9b20Kj/MScE7
ajmVVlOWefH+UA715Udp3tLoRH1Bl+nMq/jxw5UInLhBXXUNhcTJ2BJFfr5d15Pq6RarTRFIrTs4
jUxj3K0SA3f69frLzcfS7dSDPDqVeDgMfa37CI/PXzqSO5z9tJNdwCGIDTZSMxCkdJiAJLlAF/IX
iKguuthBI6/7dYzrAhJYJkMbN6wLj5PwMxly4t47MHGo2BUe7L8YDEohFZRftS0qnIVVDDKU55V4
IGOxN/uT81G/WOGzcMW8Vcia/u0dIegSycn5nwNmpNDO3HDTDMUbv8Ti0K27C/yKbYjlrA+VhJUo
AQZxIURRsGTOHpwbHGXqRE88/b3pENNzLHAlfytnwRbx32yA4kb9as0MXile3IG62+HfzoOfeRe4
LxiMdGt5rGy35SlHY5rv9EozhUIGqRK/b7EqVv4hZ/tW30dYyduam2rwKgDHUqFaJnxoTo4ENvOQ
sL7da6wUJomneTnQvIcrQq+b26KoRW5Gz/t7v4ckyLN7dT5F2S0eDLsZrLxFFBaxiEQBuBcqj5cN
N4hAx9cpxkxlT/Yr4Fysg5kxqFXP6yqKus+SAA1qqAzRO5Ka/UqflJGhA4a4rG/eeqeugg0SaglE
y+qvd+eII/mAEW+zn6CUr0R96ZIBZRgUzy2h3GO8SPRTFI3pQgIGQ7seOqavOxXy8I0SxNubU91D
YqHkR810Xkmuq9OBxHcvN9HDDiHYk0+Ezs3gqh1yWK0I3Q81Fgp9NIxBJQ7aaDjCGXScKtVi22YA
pPzUFxP5ni1KtkBL4EgqyFALVPCztIWNX6vrzmRNHKqgAtjltWlYgqdQVeEh5/Bp3FfdAttUDcLn
kdl/LBPlOBdgvK71qmwC5vE74kemarboYD7K2Vj7q13HlLQ/uZR0Q65acnRhof2pAibxW4X9N5R4
X+gj+qWXM106RHfno2rwwz0LxP2b8Q+Uba6lduII5gGtwWAXJQ2Ob6NzBSBoWPnW+AjJB5BHLr/q
W2j1X5z1E2NIKWmkgkYjbZW5dsrkqSTRoK1K+L3bebE5D1Puhzspm+zjnEJ7C+Jc6D0ufyeyqnO5
S438jQ/cwCfArJBWvtl4cC8oq5zJzx+ZbkVOdqvWa3LfmgDc5xS9nWqM6rXkGog9hKXfofnk9qX8
hpsYnOLxm7d7FnFf7dL3FoOQ7BFU/W3WFiGEmd+0c4AbtLE+HvR9ZS87dHvk3Trv6fQBiVWyLDVP
ZPytott/rvDd2gVtl1LZIDfxytE1Vr+Ih6hIHALP/OyguUu2gnt1VH0ocKtexgc0xxUUTACf3Ajr
AJrK5VnOKj4mK8KGOSTZNURKLel/DQfzVyNEC5CceR6cOqCRphc+NuQVFw2mgwdPqhrun2GvCCvJ
OR+b7zvAN4iemq0zPSgFu9VANCyum5RWZ5M+3BP5/0Ki+7Akv0f1eQWFqGjVlKGTt5toiYNwhGsI
IO40VMZME3vVvvuVhRHDlPjZBYRDeZzklPESrBsJNEYYcaSGvD4icc2SrBGxXhvjjyVF8O+p8/RK
j4vQFbMEnI7hkYJGV6MGR7MqDeFl8ljBKAR0HFJWb3uJ0M7tM90BtNsgWL6FZQk7ncp3QqYBxQOk
lRcZGiLTmydWUdnoL7KqSGUEGYXDCPISlpgEWerT/XfHmxBofn1s9FqY1xIswQyuCdOqEZ+Bzn4V
wsARzbDZ6ldFKkbMPOMv1Op7qB07iWyDTF0qpjnCK2n7H6e7HeML0eMh9GYekPNhyD+FCTKxPEua
3PcoJ07/pXY+WgkARP1tgxNRfJs8jDzcOgUxglKbw2JSuXx0q2gtWzzjCuvZ2c4GGhhgbfR8rkQZ
ETez0c25SDpGJQpQvZ09YRNQpnB+e575sQodIZloBDoyXGcCclcVpSa00hD3NVPZJu8y2ggbTVDW
eF1BsR3L5gWTp22EX37lLKeAF3vmcs1MR4zxTVIAcFLLzmLBxVebdNKxzdIFOIhHnsRfdfs7vuc1
uOadJQUs9V1sM/yc+CI+LpK4jq2mLI9r40YBDt5oEOQirxAhkeUMcQ7wvoXeR1+sUKiprhAoCfnC
2ZxdzCR1UMIEaYQFd1tH/qC2NPqP10Zmro4pC6DMMibHiysKquOAxYeY9vSlq1ELp9CibHQCZusU
5tNUK+lh3iuhdh51o6uW9ABN6NcB0aiKFyjC5I+msrShsc4/k+waDL1/EXYTWfDGb/Pl5r+eVEMo
klLmSlYNmCirNdQRrT5fAoGhl0z6OdpsI57HeWQEmpLQgsnrXX0oRGu83p5JQWfTel6GB7ocmEgH
c7x4uNB391vtOAFOOgsQBI0JYZZ/znVmmL8r4hMzijCnXLv9RNeGPouCxWL+wQYne4Kb+pdC7iKi
/WeSvonPAs/RVOg3YRrIIVlTBEgC4sxCEas2xhf3MEIDCXrqep9/T3dJLyMnDSRnIBgvZ5Y24cHS
1flbcpxcK+dUJ4M0rncT/xN2x2qJaiId5OVq8afFOEoHOP164wfl64pG5Iy1M1VpNhpng0+coy1w
mXr0q84oQG0IX+Nbuufq+TzR20HW4atm37vMnJmwUmhRUhSEZRxRUWHpkyn43x2WERP1lHHZDLVa
45NM8ZtP/8ZMsZdS1UUEcYe4lewr7oP3GirB6G/nD9tJkq/yLLw50cJ2OcGxKW48n1Ah67QimcI0
X+gWraOXMCUpMVsz3Egk4EskOHZT19G9tZ7U0kmDszIiCV5wduI0OJ1UwF9wOJ/ZhR4+xD/N59yZ
TfSbnA5iSG6iKihhEWociGJeDcd2vvi4hVQjyZRBSeiFd8B/9qaaSkO0yMesb6kSg7wl3mfwWVYM
QhNbcR3KeX7Z0HgO8CheezTDekwEmPi/Ww4jheKU9+nVGuR3AE9JdlrjYUIJuUcXGYOrYkVMCu/1
mjg81Rl+N8Q37xqQ9OZWjKZ1FrZt/5qNnC6ux9g4fyQX5hYekQi3+sRoDnpMYhmShvK/KwryfC5O
McNOtxhn77lnrLO36kzjxP2V5W7acIgS/770IZ5vbyTJYeFpayQcegu6g/ajiDgnA8KOac8hpcFk
JxOR2cfLppPofhbpk/59di4w8eUuYXRLP7hOJcjW9c622j48eLcMPsfgdrgHBsKuVXBhp/9Ytnp/
A46bHPOAV06eq9X4kLpQgssihuApH48PAkCW/rPef8rwmkNq6g0IQVioXHNg9jHs8QUcGIJwpDet
vUaCOM1FggckQNjg+6YhSJRRy61DfqZW1+cT62p+qeaxP4dt6On1s5HQk5wPlCOPEfKL8AOcZkBU
w3h+Jpb9wZCar20BFrLdx8uQtIr9EEDQgN3iumzfN5OdBjWDh+ekMbgG0gHwU5Xh7zx13eESrff4
d4wR0USkYefxLQIXrgaC/XHULq81HN6qbDwLeXFFG3WnxtdmzyD7xaxRiNu895JoaLDCUR8oTGWC
eUypmwMDsGyllMzeWF2O3gna6iin6//fFLL0Nx2F5f4031efql4TkYoZwkdMYjlpvVnPWiMjj+aD
mUCoSdOBSCn42afheaVs60TxUDagwDrKE5930WtNCBUltheilIVAc9NY4jW59vvqn3XXYn+uWY7S
fV0CpPF8LAWSgxSCLP/ZjLcGU5PXNec3Itqa1BsxPh5A+m0yx8Lnv7yYtVJciKZrbit5sj+B7Fm2
w3jA55QTwA6keMuam4pRlp2X0qk4i029Fq2p25jHsHXJjx4+gtr6x1KvMfU8jtiLCbpCPMakW7lv
RnYVt62m/lf6Z/K4lrozgTUC67EsPCrw3yTaQ+/FhAioW+Gfovr9QLEh4YzzfX0WIhltOORswMcw
5BSrrGKRoBTtJ+3lci1skDRD8DQQveKIz1mCgs2OcxorwnsxJkbXqrkwFowko71MXDveLugzvtrY
GPPPnBGuKVXzqPGQ96A7Ow8PU0Djacg320OPzIc2evjygUxQu3XRAzCiI0TbS2eHmIxzwS1luxbO
7tnuL6LQgnoADO3BwtW+XBvkvkwnQmhaTd/BlpdHH0QbGQUSY4WU6wrn95f++UhJCOMWHcoM++Uv
U7g3tyQV15Ss5pH/mINlmQdl+1Gr0LWesCr7LbPItUXfVBWuuMWfyE6BuHQwp5bLrA5LjXKCCe9C
IF0LmYB4cG71T5BXAa8ARWirD+J0ilP8YdmvC1iaNKnDcZHM5YtdI8o/cQZbtInehnedHerCORR6
NOLyq1efHldJTo5oQicGvHWkL1HUFNhAw45wkV5Ws41jMO4REabeJFDl/XvUbHpj+JJV9PZlwefn
uwMx955GEQJ04mgNllK5LFhOWJXlINLQWbuA+7+MIuVbPJeRSY335U57eX5LioZGZBH42QCRWgx0
SFWFM1JYWYE5fIsUXZ0iL3GH8XzXtUs+35GhXxzuHVQlYMyn0tMGA8EtCCtRXH2qU2zMRnU1xmfZ
ceYsnTogpCoJT8zDCdSFamFRpWeOztNkKjKohVle3zkBPwIajHvsr9B+pCD+jHsm/H94Co6IOIeF
c46lTWzpdZsG/Ch+CKAkUGVi/bULFex3hhLlppJOQUgcSYxkk8rhws3CdUNdQ0pNORYMBeA88jW4
vSDPFyupcWoZ7kf3J1bTAaPGxSm6AY53VLNcj/oiiKi8vntdRs0QciA4ahaz9YSeaHRb0ELJS/Zp
dh9iEn0sykg5kHX2nseRYAQNsCZ2TpREABLX9WkedatoCnzLhYbYO14RYqOzrmoseMb8RdaMovFC
uA/zy7/z10Fzm9LxxwZ1sqOllI5buYCXhR8IRJrFsTaB2cfq4lDBQLGSZX/Mv9D5X1qcwBqyleN6
Tjogq9KGXUfnDyaqRlEJvqkoZD1tTBbW1RkcHQesvok37ftvZCU8osJbWnk7BPLOvuN9Cd48/TjK
D6ofRd+/OD7i2RCw6/E88mjpBdTA/+jAnqm86xX2rKzD636rHgnDIog2UtXzbGky0lonBiP5F8sA
vAZG5otiCkheTAISfvoSwr2c2I74jVBgRdEZZaOVtoS/TMy2nbdqoIU64V509NUzR8aNEBTYUz7i
rmQz5MTRZEVGtsCejxSn8GUbPvQAZUHCA7edbLHFGXbmAFJ2HKEFSbFfTxg5gOXJeOsolLdFRyT5
EXSg5hJryi03/TRUkh2PTJc6SEG6RMr/48yvOsPFZHs2UU8+OUiejRM7EpF4UIVJ3DvhMVv1//6g
82yGsF0W/6iM9is+FgsBqoQB7fyEFjSQPgjwFhRGQgTVFrpdkzATx32QK1EGgAqUfLFT4wkQnodB
IrTNduWC2MCGzZL3WCXOhmfBhIYPwbQDYPzGpy8meU6StiYl+R8Q05NF01j6IQMMOiKgeqeobQI0
W+vjriNWOoTVv9o5tkwqsswzpV4BLBDga3VAbl6ynM3KEERV8eGRiDpLof5t0/ML4yR8vzCFjYNU
62AhPF6TEfaODe5zNAlowRE8A2rXLcC5tBAlj8JfhqjTDgjCp60Eu/++k06/DonLJDGLr6pa5aPC
HaXZuHeHGzOWOx3l3ixknGjyev+Z7o576zLVr4ZFWoPVh6JCp9EieKKBMg1I8dbHGHN8vCq/99Cu
X9zJ/6E+dCd+5DgyuF14YFEcwmSR+Mvw1r65aNmmFk4yODb+M+LWs3hTJrf6zmQx4sseuu003UAx
ZoYbonn3glOLcQCAiPGOtPXz91MLfgdCZAdaUk6iPleneigWijF9E1PED801vPcfBJUBXeAGB9kU
Czs2+gX1ph9kx9zdKqxyFK8SycrjOOs/UKy7x9PD84NTiZbwGwMbYM1drO+eg1aCCU+4gq5XEcmE
igabHljzRtviPnzj/IyRlDxFhBS6J47K6SFJGVzyQAw+/HkRxJCpoUhy+KndhWLRoUs/Y+9HyVre
1FjUaYnOesHndPbe2DIKysONqnOQJFiss7uZrKT1BBHyFs2LlYMsZpn06Ckmk2qwPmgK1PX2K914
jNz2SdDpaErONrPu3wHVg2NYcH8tNqCDah7r/ZzapLC34EKtstAnCUipQG/K8j7GWdMEuzuXwX9n
EKvt15uKLljWI6wUMtndAKLuIra1pDsrLcFfd30IjpJIxMxBtQfk/OatfKDldOeFBP4TOD0EIlHP
Q6J1/KekO5VViVAGZVTtRQtWsDO+NJVu7ynA+pcZK1saPMApkdy2WbY4NBR0GjfwVZEKbDrq48GN
v2NlvjJjmlARy6b9UK20zGSEETgZvmavWRPOSzbdAQ7DiQ7fzRRDX9J2oKqd/zMglMpZ89L8rYhC
py++Z/6zoSvKIZFHtfM0bBGjz24v8XmNfyzLjavV36/zCD5WyO7VprfBBWRDIP16Jq4dp65yIcqI
6En9Cv1TQR5GtzhoS/yV1K7sxZjtgrx4trI8AuPTuKUeuA58CSqXbRKNEz9tyzBtUvYHdnfmzgbX
YGPSs8Puts3yHL/o2S7NV2eTkDxxJYC7uUewSYT9jLvKhpyY81p30/PDZx3PJDolbXDt8RRUpuyM
0pHcJm0xiKS4Bbn5oSfuhrWU5qqRC8zeplBph7H0+jMg13p222lwpD6oMb1X4AImWzD5h7lj4tV2
VcZCi6yGw7T857tC/DvIdnr8I27zzTTTs/fvsCGlyb2JoQ8bty1JVAHMm+7NLbioTG0FkyqCjjks
MHjqn9cLxJCayJ1kYU1Fxj2ZyWebQwocp26S6F12gAVC7QXLozxotbY+ZVEsP/G8t7zhFS4Ro9og
vlggVvqTH8r1hxQzW+PgaxVwr5Ptz+YwrTaeLtHE/edk8zFK8D2tFr5HkVfB3+zIri6aJNR0YTgX
Wlg3UtCX4OmB0EF7wZ6hkxRy5/ghQZBqEemdJ5eJwjrIOu28uy+GbVdqwxcqTsyiSfRq4px6jGM+
thb65h62Lx+qzHIj0f3GfO0+KhI8o/wbmqqaiL2dSNbL3RtM5bcrbiPkKf2EjapOyNjeZhyhFV5r
YkSB/7QxmQczURmWKCEUenMQVXpmhyJz9KBk34VlXX2ZpHDDjqmONkJLmYb42vqUpyPUmDQAnaxt
kPwdkrOif9yV7RcNVEaLB2WjCn0hdLSrEe7lqAXf0WjRE4gfTnkkEqkZ0WcXvrH3NzmEw6XKcHwZ
EfEz0kxZYsviwur+WuLrA/vHkpUz7/p+Kvev2VHSxNP5ppOd8Lq4L68Y/pKb8g2AXkBf9WtDUonD
QSPzjRAkTpvJIUTAS9gHX34/EJ555kad7wqGT2Ik9gs5gL4U3I8RaH6VnvX42IGL76C5umWgjTFd
BXm1z4Ip1yeGluVn3/Khs8MPERTc6FJzmJB817ZUEiqdQCH4kmfD8IBhv5BjhRGIxr1m+8FrKseD
4Vgd5yN48l0SShhiBbu1MHenGURLS+nB3vW6EdqU2ThUwLQfCu3Ydy0XKCYhu6xEhw4VrsQBuyxx
Vp+MMp9n4Y6+81TCY+OEI28aBR6Ey6YrzssvRppvQYY9hyfRmp7Bmuz3V1awwguXroluqJRrDVw7
ClTfisWPW8gaIrdzoPjs9pbNdUDHQEDmECAVqGutfQcfv50VALn+xgLDxyIbHIGxkYQtcIXabkS/
mpkwKXvmf5kTMYXB1SSBRZCAdG4q2Gtcdh8/Y9ei9/Y52StVb2PDX2iDEqysfVIBmLMEFDKmHdIr
9liDa1U1N8ZsdJjHtxuITCB1IoRIwM0mHgYmSg3m5J7t2sSKlwg+mmf1J5MViDSk6hDM8lflqlCt
6BhjGg1EWWGdz3uqo4x5dm3+9HRQBnaayb3/Obt0SxMzEMOu5bXwv/ilnaDXDVEemv8xLBsLO0nK
h2Yt/oY3mul20uVF68tj6N1gIwBFJ0oIw1PGmEveDIwx17TUhzhuJYLM0Iuf8a5CLx76sqqzM7AJ
F9ZYvXfw22apPXxB1w3RFrQkCwN1gjt22gDcySKkRyarsLDDBQ4aBgCNoqZBVzglCEsJU51TFnxM
kh4nSuvz17zeDi8GYxPFjP2UTO3zW3by6YjYeSJSjVzoMYf/WUyl0wCBQ+/y0jotFPIXHzmtrebB
6lZqfJMGq7HryY+pEZNH4hpaf2SAHaSa0Ru0olZ+9dHNpKrVcYLz4r98nAZp9xDNNn1/MYIU/HoR
lAiTFRixSohNVxs7ZOcNd6/PKsUM9tUx2ybKWDUF4F9x28nXQEpVJM1V9rsFSoB9mvZF0msKVMkf
HUS4l9jj2WW7b1OYun0IN+BhqRR0TUxvLycWLuhnyYIz7/hA+/U8pxIdxdpJVr5nYc1bmKUoWXH9
1BVvzXSaT0VvghcJmAHKJ5/2Nb7DiIME3w1gywjId0lva3JkYF9t2dXOvGf5PgRfChV73gtPwlbK
rdKveo5Scf4d3zb8mvwveyc+JU21rg7GCNuVqtZ5VdA4aA6RlJB+mLEQt4Z1FhZZLbcSxncW6U/4
RKlEj1Rd5rxjgAvg3CKiQBdy1DiQ2WhctvDEGuCmwtrbeQqH4Eg/1HLqhR95NZLzvDwJxy5YvoFA
w+C3j8oLa5la0dsYrtaztM2NyDELf9biFko5qkbyviOQpzAj7Nh7B2rqYNbBElPYsgl2leaLV+Lr
r5qSC8Bgy20fADD7OLNrrHmNvK8+NuhgpuCkk+6LywVZsQ1Mn4T/EJuNcSD6vJwNGevq7iuE+eb5
zMuhpnBTKBd73pleWlOCe74wVW1I0CTnf3hTWR7ZOct8GyBFDSjdOV+GO4MOgx/g9sJKhdvaIbBn
rAKdRmNDUyfWl1VPnP29rdeJvk7YRpEqTNfJ3bKBCuwRj8P/fDGbrolQckVoFFWg1d89zjv27BrH
rc9hCCDaW/GT+9LAtlhs71AVBANIN47m2szhvBBF4Q/zxtRxLmFNu60WPTO9Hl8dyHTKxK80Oftm
IlzTyZ6UPtcZmFX7drSvAuvsaejhsMzLJjqvmUOtbkRX0Hv4jzdpoO2uC3h05gRPNBWvW5Asaind
8cjbyAWcO9PsNFO8I9URnAOIXQjq/dJAg5xaseKlwqDGEKjPU6vmxnbLdLnL9H0Z8fT8264HqYaa
TZ1WG0WnI3vOteuRPnTb9MH7FCvEy8BrQ7l6NHCxb5IhERkbf97CGvcPtNR8rBwKeBamUE9xPfE8
LikElrLCY22oLYE9b6RxQxHuoAiCIYnjA1N87rCJ6fjsrDZAEZeujpZxs8xp7Yo/BbQAV6KaZUYo
OLl9Hf332crOv7RRN9MnxHw74itS9UxAexY8oqyTV2ANkanyjW6ucE7pDklxHeEEx52JK2BYpaFs
Q9M/7SVhCsmJVfr4KwK2qNIKE2IRtZKCdG4WoAsxFgiOnbIkbVU5nMqVt2sc5+ooQML+LrqtH6Wj
Kdv3w8DNCLrPMyZAVfZ0O0lUO3n5qgogaDiPoUwUHEPP/XU4MTGOm5Ym7zf2fkXKxGJ47fFAwrLl
lPLhz/vE8OxZakxScDbPPWEhFBY4J6/vy0atLphG7z1yP5V6nbP2c7fzruLe+GfsDqoc6BMgRyIi
ApXOlmO4U/tDDjpXyRflrK1ydWkqmq0rtW84zmXw+b+m1tKCWsbHwVOv50PbNs3Rwd6pgqanP7SV
H2ClQjcxHQ/U/Gix/L1aTpbcVCYiQxSl69lUZ6PVIkC9lSGzL33GvMfaYEuC1kDYwhmSA8hLs3CS
Tnu8y6/SBoLdBQJiceDZl8qhyQyhjnpd+gmy4x0ymdKf6jZZZQU7K9wmlf9jzuW+f5DGdolpf1ug
iTLX3UtYn1dYEzeCyyM22sUhkaUnV6zIh2FX9S+61MPFll8QkitzKOe1zDOh7UItwCBMme50PFiJ
CDTh2/GEIRAIT4JeD1KlhJXnK7coNrDPTctqm1y+bHOFQtJJJ/JGpYCowED9RQXbqOd5vK6zOEGE
yV1gS3+qP1Mlau5hPSLREmn5H2MLmCms32zoMyX6uNgF1kfkVa0v9LT5Y56hDcqQv6oxsN5JoqGg
1Ja6b95vx0l6jtlw6OwVa/jaQj+CzjCOOhdB61vZY6+gNb+xF7gwhFFMtMAd1MsITW8Gz0LpX/CF
qx0dDWGnksczYIzJnb/aZHyGBikCA1BqrFpAmRtTEbY0RMLSkDa9vg7U1YXlWnjaBcRIqT5EZmEn
0kShK4zqmWVYFieXjyAhIJ2OJ/IeKqFq5rYvp08kACoqw6YiE2D7QWejtpp+2ryplC3RonObAmpj
gbfWrcj//6wsszWvwzqOfvvZC/NB9f9jCMbpCWAnyeBPn+tO5oqnprjfvJQ7AYdyugrdjKPQAWsm
Q4zgOz6gmEukCCazYg416eo7Ul88IlY53LUTN8rd8Flv7p1K5hNQ8cQWuSg7TCij9JPtlc/6eiWS
Rx43iWRRJ9y50LbQZo2uYbRBZsHDFygqowvCsSj7wJbpib9Mr0PESJfyOGTO+E37u3qrNddr7HCv
hm9UT1eqhNGNUBgboQgWP4OQRSYteH96DuyUgYaV08UoND6RqfDOuIU+fYm1N+/WPwATgpskwvhy
1a6rnO6Mdnx9PgdLqIz319hRduwzCA4ymZNictrv7SLP6xLM17BlTf/gnzFFHDIX/bfcfdM+Fqqu
Vnh9VBo7fhGZNgYYAE5Dmt60Qd3OoXiOIrd9aW+r/jUUuTQ7jSQGKNE+9gNOczIZI7U9jKCRBnMe
zcwOEXWwZ2BAr5W8Wph5x1LdhrS1TU3QzQrnKQ6K7QLhmRXjzqwAkw1LmCQykxi+3Xj+s1OdKPyE
BWovSZs0Bjfp3HzhAoX1naH+0luYqZ/CBkP3RNVAKXr42U5aWYmQiBjLZsrU6FrghW0HUX3L3BS2
48aCq7sQN6aTFa3dXboGgRV2GZ7DNKk2/7dQhKTbXv5f2dUwtTeBP3qiFBIDUPQVH/qLHFOqyJq3
g0W0HD8UrYMu6H/J1JThUs5KWTvJtX+BREz0EkVLciyUwncXkIvH5IH1FCTnQ1Sa3246gWr3d/uw
3RvIQLY+D5kZqQXSG/2h7eMF5gbz/oWuUgcfprey7zBD037sUHKVJ2yFqbIZn3Fi935YhxLbO587
D0X7jFKFb6rOFioGlpVi2+s03+kRy7AAtgOkNlEqUIqtNkRrQowCIKVtG4mF7KxzzHA09ZLnYkfp
3eYXeDWVhLb7CYC+6VPPUV/aIDPp40vnbubDIpPp6dTcBzViojmXDLOHK1co5ZOAk4OjIGWJgf6d
goCQCc4QjiOxs5srcd2rwGzj6iRUBOcDeg6z3RrqgQZsNivsGF8fRu6bsTjEk/KrW9G50PCBpBkQ
Al3S3tAIkJjvRooBh8Xp3pxe81MrCcFVdisHT3swPdAmqe+c5XoxfDEymRXf1bO+GCAyqnM6Vpm8
7l9RXG6efkeNvIx98Hj4r302rKps8LU2iyx5e2aHT7+rbeveSgZWx7XEZMsoyn3NdvjRLoJ3UAX+
NVe8gaFouGOOwymvrzZQST4EPM7iegk40bNqxRSwUMmDXbY8K1rE6cXs6E/it9GL0a5DSuBxAygt
YajK92ql0P/WC2L7CeWMjzF6IdfVNHO25rROHIFHMmuAZ5ep2AC+ZkUMxlN2tBwDwQWwTDYSppVh
C75DfS3mAL6YAf9f5BarDEdGlBXHFenNXs1jNyilrIHdtQOimNu+vn0YZh1bRUDfxWPR+hPOMiD3
VTxw9ucLn/MqdEDMTP4wH+OGFpl8hFN26EPYMYjvXInNSNneAp3UsAArSFnyjItE6S5Vj1Ex0d/r
sDWAF1LNVAabMLnVfs2Xhj71c9GQNSR//faig3326GhpycR39cGRqRQ+dM7W8kdNzqI43b5WH9J+
6DPf14b3q8eyyu3ElGOgkngDglIQ5JcAVIXSSpGVK0iOan4v5ge5ATrdCJpPF3j8w6vnERpdLLsl
XVTJ2ntJMBjNAe0FqPMvU9uCjHEyGaZ3gVew8MotQqeKCdNDiDNDbIuGs66Bt3l7pt+CKnCR5lzf
ank/hK4AW06SwJounws20xJ4WiYVfzEgDbA4xGHTn4x2WivITjAGwyw9HUVTwc3E8Rle5BKCnODK
3m4YgjvMmU1D+2HQsRASlnqGjW5i9OqCdszXYymrHZh2JtrfieapRCDvOLORAmqOmg3+ZcjxRWrN
fe4eoP5dQxZLE13AxdrpmhozGjl9S1HTVqQJyt//0odW75Vnn+P6JjBbGrupsP99BaYyWT2zFJke
WPkNDhkJJlwGUJFB/yPNTpJDZiXggLk0lFGznDZXJDKtXJrjzFdHkJRDlqGD1Syki6WZWBfdDx8x
gUmqkJHcPXC6oqSUHh8nvfRdAAGVDhvlzsTJrE+FqSOAAKS76+merDvn9r+i0hyE5dKM/ZaSkfnE
L4d90VP6BifbahjwH6DWz+eQ7XuozYnt9Ab/gkxoe25DC8jjxekc6bPOXD8a/yAcKDr617iVSd8o
v3iJBR6AjGik22m7Oytwsqy5GU6wYjIsUlOPoBR8jRgMFxMPUmPR+kNUkB4dNqwiEFyKybHD/caM
BsucF5NbWimlDKH04rxWUvSj+g3QOljvdEfHuheV3ur13FFdVgchrdeP4w==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library synplify;
use synplify.components.all;
library gw1ns;
use gw1ns.components.all;

entity Gowin_EMPU_Top is
port(
  sys_clk :  in std_logic;
  rtc_src_clk :  in std_logic;
  gpio :  inout std_logic_vector(15 downto 0);
  user_int_0 :  in std_logic;
  user_int_1 :  in std_logic;
  user_int_2 :  in std_logic;
  reset_n :  in std_logic);
end Gowin_EMPU_Top;
architecture beh of Gowin_EMPU_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~Gowin_EMPU.Gowin_EMPU_Top\
port(
  reset_n: in std_logic;
  sys_clk: in std_logic;
  rtc_src_clk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  user_int_0: in std_logic;
  user_int_1: in std_logic;
  user_int_2: in std_logic;
  gpio : inout std_logic_vector(15 downto 0));
end component;
begin
GND_s5: GND
port map (
  G => GND_0);
VCC_s6: VCC
port map (
  V => VCC_0);
Gowin_EMPU_inst: \~Gowin_EMPU.Gowin_EMPU_Top\
port map(
  reset_n => reset_n,
  sys_clk => sys_clk,
  rtc_src_clk => rtc_src_clk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  user_int_0 => user_int_0,
  user_int_1 => user_int_1,
  user_int_2 => user_int_2,
  gpio(15 downto 0) => gpio(15 downto 0));
end beh;
